`default_nettype none

module coll_table(
    input wire [8:0] in,
    output reg [7:0] out
);

always @(*) begin
    case(in)
        9'b0_00_0_00_00_0: out = 8'b1_00_1_00_01;
        9'b0_00_0_00_00_1: out = 8'b1_00_1_00_01;
        9'b0_00_0_00_01_0: out = 8'b1_00_0_00_10;
        9'b0_00_0_00_01_1: out = 8'b1_00_0_00_10;
        9'b0_00_0_00_10_0: out = 8'b1_00_0_00_01;
        9'b0_00_0_00_10_1: out = 8'b1_00_0_00_01;
        9'b0_00_0_00_11_0: out = 8'b0_00_0_00_01;
        9'b0_00_0_00_11_1: out = 8'b0_00_0_00_01;
        9'b0_00_0_01_00_0: out = 8'b1_01_1_00_10;
        9'b0_00_0_01_00_1: out = 8'b1_01_1_00_10;
        9'b0_00_0_01_01_0: out = 8'b1_01_0_00_10;
        9'b0_00_0_01_01_1: out = 8'b1_01_0_00_10;
        9'b0_00_0_01_10_0: out = 8'b0_00_0_01_01;
        9'b0_00_0_01_10_1: out = 8'b0_00_0_01_01;
        9'b0_00_0_01_11_0: out = 8'b0_00_0_01_00;
        9'b0_00_0_01_11_1: out = 8'b0_00_0_01_00;
        9'b0_00_0_10_00_0: out = 8'b1_10_1_00_10;
        9'b0_00_0_10_00_1: out = 8'b1_10_1_00_10;
        9'b0_00_0_10_01_0: out = 8'b1_10_0_00_10;
        9'b0_00_0_10_01_1: out = 8'b1_01_0_01_10;
        9'b0_00_0_10_10_0: out = 8'b0_00_0_10_01;
        9'b0_00_0_10_10_1: out = 8'b0_00_0_10_01;
        9'b0_00_0_10_11_0: out = 8'b0_00_0_10_00;
        9'b0_00_0_10_11_1: out = 8'b0_00_0_10_00;
        9'b0_00_0_11_00_0: out = 8'b1_11_1_00_10;
        9'b0_00_0_11_00_1: out = 8'b1_11_1_00_10;
        9'b0_00_0_11_01_0: out = 8'b1_11_0_00_10;
        9'b0_00_0_11_01_1: out = 8'b1_10_0_01_10;
        9'b0_00_0_11_10_0: out = 8'b0_00_0_11_01;
        9'b0_00_0_11_10_1: out = 8'b0_00_0_11_01;
        9'b0_00_0_11_11_0: out = 8'b0_00_0_11_00;
        9'b0_00_0_11_11_1: out = 8'b0_00_0_11_00;
        9'b0_00_1_00_00_0: out = 8'b0_00_1_00_01;
        9'b0_00_1_00_00_1: out = 8'b0_00_1_00_01;
        9'b0_00_1_00_01_0: out = 8'b1_00_1_00_01;
        9'b0_00_1_00_01_1: out = 8'b1_00_1_00_01;
        9'b0_00_1_00_10_0: out = 8'b1_00_1_00_10;
        9'b0_00_1_00_10_1: out = 8'b1_00_1_00_10;
        9'b0_00_1_00_11_0: out = 8'b1_00_0_00_01;
        9'b0_00_1_00_11_1: out = 8'b1_00_0_00_01;
        9'b0_00_1_01_00_0: out = 8'b0_00_1_01_00;
        9'b0_00_1_01_00_1: out = 8'b0_00_1_01_00;
        9'b0_00_1_01_01_0: out = 8'b0_00_1_01_01;
        9'b0_00_1_01_01_1: out = 8'b0_00_1_01_01;
        9'b0_00_1_01_10_0: out = 8'b1_01_1_00_10;
        9'b0_00_1_01_10_1: out = 8'b1_01_1_00_10;
        9'b0_00_1_01_11_0: out = 8'b1_01_0_00_10;
        9'b0_00_1_01_11_1: out = 8'b1_01_0_00_10;
        9'b0_00_1_10_00_0: out = 8'b0_00_1_10_00;
        9'b0_00_1_10_00_1: out = 8'b0_00_1_10_00;
        9'b0_00_1_10_01_0: out = 8'b0_00_1_10_01;
        9'b0_00_1_10_01_1: out = 8'b0_00_1_10_01;
        9'b0_00_1_10_10_0: out = 8'b1_10_1_00_10;
        9'b0_00_1_10_10_1: out = 8'b1_01_1_01_10;
        9'b0_00_1_10_11_0: out = 8'b1_10_0_00_10;
        9'b0_00_1_10_11_1: out = 8'b1_10_0_00_10;
        9'b0_00_1_11_00_0: out = 8'b0_00_1_11_00;
        9'b0_00_1_11_00_1: out = 8'b0_00_1_11_00;
        9'b0_00_1_11_01_0: out = 8'b0_00_1_11_01;
        9'b0_00_1_11_01_1: out = 8'b0_00_1_11_01;
        9'b0_00_1_11_10_0: out = 8'b1_11_1_00_10;
        9'b0_00_1_11_10_1: out = 8'b1_10_1_01_10;
        9'b0_00_1_11_11_0: out = 8'b1_11_0_00_10;
        9'b0_00_1_11_11_1: out = 8'b1_11_0_00_10;
        9'b0_01_0_00_00_0: out = 8'b1_01_1_00_10;
        9'b0_01_0_00_00_1: out = 8'b1_00_1_01_10;
        9'b0_01_0_00_01_0: out = 8'b1_01_1_00_10;
        9'b0_01_0_00_01_1: out = 8'b1_01_1_00_10;
        9'b0_01_0_00_10_0: out = 8'b1_00_0_01_10;
        9'b0_01_0_00_10_1: out = 8'b1_00_0_01_10;
        9'b0_01_0_00_11_0: out = 8'b0_00_0_01_01;
        9'b0_01_0_00_11_1: out = 8'b0_00_0_01_01;
        9'b0_01_0_01_00_0: out = 8'b1_10_1_00_11;
        9'b0_01_0_01_00_1: out = 8'b1_01_1_01_11;
        9'b0_01_0_01_01_0: out = 8'b1_10_0_00_11;
        9'b0_01_0_01_01_1: out = 8'b1_10_0_00_11;
        9'b0_01_0_01_10_0: out = 8'b1_00_0_10_01;
        9'b0_01_0_01_10_1: out = 8'b1_00_0_10_01;
        9'b0_01_0_01_11_0: out = 8'b0_01_0_01_01;
        9'b0_01_0_01_11_1: out = 8'b0_00_0_10_01;
        9'b0_01_0_10_00_0: out = 8'b1_11_1_00_11;
        9'b0_01_0_10_00_1: out = 8'b1_11_1_00_11;
        9'b0_01_0_10_01_0: out = 8'b1_11_0_00_11;
        9'b0_01_0_10_01_1: out = 8'b1_11_0_00_11;
        9'b0_01_0_10_10_0: out = 8'b1_00_0_11_01;
        9'b0_01_0_10_10_1: out = 8'b1_00_0_11_01;
        9'b0_01_0_10_11_0: out = 8'b0_01_0_10_01;
        9'b0_01_0_10_11_1: out = 8'b0_00_0_11_01;
        9'b0_01_0_11_00_0: out = 8'bx_xx_x_xx_xx;
        9'b0_01_0_11_00_1: out = 8'bx_xx_x_xx_xx;
        9'b0_01_0_11_01_0: out = 8'bx_xx_x_xx_xx;
        9'b0_01_0_11_01_1: out = 8'bx_xx_x_xx_xx;
        9'b0_01_0_11_10_0: out = 8'bx_xx_x_xx_xx;
        9'b0_01_0_11_10_1: out = 8'bx_xx_x_xx_xx;
        9'b0_01_0_11_11_0: out = 8'bx_xx_x_xx_xx;
        9'b0_01_0_11_11_1: out = 8'bx_xx_x_xx_xx;
        9'b0_01_1_00_00_0: out = 8'b0_00_1_01_01;
        9'b0_01_1_00_00_1: out = 8'b0_00_1_01_01;
        9'b0_01_1_00_01_0: out = 8'b1_00_1_01_10;
        9'b0_01_1_00_01_1: out = 8'b1_00_1_01_10;
        9'b0_01_1_00_10_0: out = 8'b1_01_0_00_10;
        9'b0_01_1_00_10_1: out = 8'b1_01_0_00_10;
        9'b0_01_1_00_11_0: out = 8'b1_01_0_00_10;
        9'b0_01_1_00_11_1: out = 8'b1_00_0_01_10;
        9'b0_01_1_01_00_0: out = 8'b0_01_1_01_01;
        9'b0_01_1_01_00_1: out = 8'b0_00_1_10_01;
        9'b0_01_1_01_01_0: out = 8'b1_00_1_10_01;
        9'b0_01_1_01_01_1: out = 8'b1_00_1_10_01;
        9'b0_01_1_01_10_0: out = 8'b1_10_1_00_11;
        9'b0_01_1_01_10_1: out = 8'b1_10_1_00_11;
        9'b0_01_1_01_11_0: out = 8'b1_10_0_00_11;
        9'b0_01_1_01_11_1: out = 8'b1_01_0_01_11;
        9'b0_01_1_10_00_0: out = 8'b0_01_1_10_01;
        9'b0_01_1_10_00_1: out = 8'b0_00_1_11_01;
        9'b0_01_1_10_01_0: out = 8'b1_00_1_11_01;
        9'b0_01_1_10_01_1: out = 8'b1_00_1_11_01;
        9'b0_01_1_10_10_0: out = 8'b1_11_1_00_11;
        9'b0_01_1_10_10_1: out = 8'b1_11_1_00_11;
        9'b0_01_1_10_11_0: out = 8'b1_11_0_00_11;
        9'b0_01_1_10_11_1: out = 8'b1_11_0_00_11;
        9'b0_01_1_11_00_0: out = 8'bx_xx_x_xx_xx;
        9'b0_01_1_11_00_1: out = 8'bx_xx_x_xx_xx;
        9'b0_01_1_11_01_0: out = 8'bx_xx_x_xx_xx;
        9'b0_01_1_11_01_1: out = 8'bx_xx_x_xx_xx;
        9'b0_01_1_11_10_0: out = 8'bx_xx_x_xx_xx;
        9'b0_01_1_11_10_1: out = 8'bx_xx_x_xx_xx;
        9'b0_01_1_11_11_0: out = 8'bx_xx_x_xx_xx;
        9'b0_01_1_11_11_1: out = 8'bx_xx_x_xx_xx;
        9'b0_10_0_00_00_0: out = 8'b1_01_1_01_11;
        9'b0_10_0_00_00_1: out = 8'b1_00_1_10_11;
        9'b0_10_0_00_01_0: out = 8'b1_10_1_00_11;
        9'b0_10_0_00_01_1: out = 8'b1_10_1_00_11;
        9'b0_10_0_00_10_0: out = 8'b1_01_0_01_10;
        9'b0_10_0_00_10_1: out = 8'b1_00_0_10_10;
        9'b0_10_0_00_11_0: out = 8'b0_00_0_10_01;
        9'b0_10_0_00_11_1: out = 8'b0_00_0_10_01;
        9'b0_10_0_01_00_0: out = 8'b1_11_1_00_11;
        9'b0_10_0_01_00_1: out = 8'b1_10_1_01_11;
        9'b0_10_0_01_01_0: out = 8'b1_11_0_00_11;
        9'b0_10_0_01_01_1: out = 8'b1_11_0_00_11;
        9'b0_10_0_01_10_0: out = 8'b1_00_0_11_10;
        9'b0_10_0_01_10_1: out = 8'b1_00_0_11_10;
        9'b0_10_0_01_11_0: out = 8'b0_00_0_11_01;
        9'b0_10_0_01_11_1: out = 8'b0_00_0_11_01;
        9'b0_10_0_10_00_0: out = 8'bx_xx_x_xx_xx;
        9'b0_10_0_10_00_1: out = 8'bx_xx_x_xx_xx;
        9'b0_10_0_10_01_0: out = 8'bx_xx_x_xx_xx;
        9'b0_10_0_10_01_1: out = 8'bx_xx_x_xx_xx;
        9'b0_10_0_10_10_0: out = 8'bx_xx_x_xx_xx;
        9'b0_10_0_10_10_1: out = 8'bx_xx_x_xx_xx;
        9'b0_10_0_10_11_0: out = 8'bx_xx_x_xx_xx;
        9'b0_10_0_10_11_1: out = 8'bx_xx_x_xx_xx;
        9'b0_10_0_11_00_0: out = 8'bx_xx_x_xx_xx;
        9'b0_10_0_11_00_1: out = 8'bx_xx_x_xx_xx;
        9'b0_10_0_11_01_0: out = 8'bx_xx_x_xx_xx;
        9'b0_10_0_11_01_1: out = 8'bx_xx_x_xx_xx;
        9'b0_10_0_11_10_0: out = 8'bx_xx_x_xx_xx;
        9'b0_10_0_11_10_1: out = 8'bx_xx_x_xx_xx;
        9'b0_10_0_11_11_0: out = 8'bx_xx_x_xx_xx;
        9'b0_10_0_11_11_1: out = 8'bx_xx_x_xx_xx;
        9'b0_10_1_00_00_0: out = 8'b0_00_1_10_01;
        9'b0_10_1_00_00_1: out = 8'b0_00_1_10_01;
        9'b0_10_1_00_01_0: out = 8'b1_01_1_01_10;
        9'b0_10_1_00_01_1: out = 8'b1_00_1_10_10;
        9'b0_10_1_00_10_0: out = 8'b1_10_0_00_11;
        9'b0_10_1_00_10_1: out = 8'b1_10_0_00_11;
        9'b0_10_1_00_11_0: out = 8'b1_01_0_01_11;
        9'b0_10_1_00_11_1: out = 8'b1_00_0_10_11;
        9'b0_10_1_01_00_0: out = 8'b0_00_1_11_01;
        9'b0_10_1_01_00_1: out = 8'b0_00_1_11_01;
        9'b0_10_1_01_01_0: out = 8'b1_00_1_11_10;
        9'b0_10_1_01_01_1: out = 8'b1_00_1_11_10;
        9'b0_10_1_01_10_0: out = 8'b1_11_1_00_11;
        9'b0_10_1_01_10_1: out = 8'b1_11_1_00_11;
        9'b0_10_1_01_11_0: out = 8'b1_11_0_00_11;
        9'b0_10_1_01_11_1: out = 8'b1_10_0_01_11;
        9'b0_10_1_10_00_0: out = 8'bx_xx_x_xx_xx;
        9'b0_10_1_10_00_1: out = 8'bx_xx_x_xx_xx;
        9'b0_10_1_10_01_0: out = 8'bx_xx_x_xx_xx;
        9'b0_10_1_10_01_1: out = 8'bx_xx_x_xx_xx;
        9'b0_10_1_10_10_0: out = 8'bx_xx_x_xx_xx;
        9'b0_10_1_10_10_1: out = 8'bx_xx_x_xx_xx;
        9'b0_10_1_10_11_0: out = 8'bx_xx_x_xx_xx;
        9'b0_10_1_10_11_1: out = 8'bx_xx_x_xx_xx;
        9'b0_10_1_11_00_0: out = 8'bx_xx_x_xx_xx;
        9'b0_10_1_11_00_1: out = 8'bx_xx_x_xx_xx;
        9'b0_10_1_11_01_0: out = 8'bx_xx_x_xx_xx;
        9'b0_10_1_11_01_1: out = 8'bx_xx_x_xx_xx;
        9'b0_10_1_11_10_0: out = 8'bx_xx_x_xx_xx;
        9'b0_10_1_11_10_1: out = 8'bx_xx_x_xx_xx;
        9'b0_10_1_11_11_0: out = 8'bx_xx_x_xx_xx;
        9'b0_10_1_11_11_1: out = 8'bx_xx_x_xx_xx;
        9'b0_11_0_00_00_0: out = 8'b1_10_1_01_11;
        9'b0_11_0_00_00_1: out = 8'b1_01_1_10_11;
        9'b0_11_0_00_01_0: out = 8'b1_11_1_00_11;
        9'b0_11_0_00_01_1: out = 8'b1_11_1_00_11;
        9'b0_11_0_00_10_0: out = 8'b1_01_0_10_11;
        9'b0_11_0_00_10_1: out = 8'b1_00_0_11_11;
        9'b0_11_0_00_11_0: out = 8'b0_00_0_11_10;
        9'b0_11_0_00_11_1: out = 8'b0_00_0_11_10;
        9'b0_11_0_01_00_0: out = 8'bx_xx_x_xx_xx;
        9'b0_11_0_01_00_1: out = 8'bx_xx_x_xx_xx;
        9'b0_11_0_01_01_0: out = 8'bx_xx_x_xx_xx;
        9'b0_11_0_01_01_1: out = 8'bx_xx_x_xx_xx;
        9'b0_11_0_01_10_0: out = 8'bx_xx_x_xx_xx;
        9'b0_11_0_01_10_1: out = 8'bx_xx_x_xx_xx;
        9'b0_11_0_01_11_0: out = 8'bx_xx_x_xx_xx;
        9'b0_11_0_01_11_1: out = 8'bx_xx_x_xx_xx;
        9'b0_11_0_10_00_0: out = 8'bx_xx_x_xx_xx;
        9'b0_11_0_10_00_1: out = 8'bx_xx_x_xx_xx;
        9'b0_11_0_10_01_0: out = 8'bx_xx_x_xx_xx;
        9'b0_11_0_10_01_1: out = 8'bx_xx_x_xx_xx;
        9'b0_11_0_10_10_0: out = 8'bx_xx_x_xx_xx;
        9'b0_11_0_10_10_1: out = 8'bx_xx_x_xx_xx;
        9'b0_11_0_10_11_0: out = 8'bx_xx_x_xx_xx;
        9'b0_11_0_10_11_1: out = 8'bx_xx_x_xx_xx;
        9'b0_11_0_11_00_0: out = 8'bx_xx_x_xx_xx;
        9'b0_11_0_11_00_1: out = 8'bx_xx_x_xx_xx;
        9'b0_11_0_11_01_0: out = 8'bx_xx_x_xx_xx;
        9'b0_11_0_11_01_1: out = 8'bx_xx_x_xx_xx;
        9'b0_11_0_11_10_0: out = 8'bx_xx_x_xx_xx;
        9'b0_11_0_11_10_1: out = 8'bx_xx_x_xx_xx;
        9'b0_11_0_11_11_0: out = 8'bx_xx_x_xx_xx;
        9'b0_11_0_11_11_1: out = 8'bx_xx_x_xx_xx;
        9'b0_11_1_00_00_0: out = 8'b0_00_1_11_10;
        9'b0_11_1_00_00_1: out = 8'b0_00_1_11_10;
        9'b0_11_1_00_01_0: out = 8'b1_01_1_10_11;
        9'b0_11_1_00_01_1: out = 8'b1_00_1_11_11;
        9'b0_11_1_00_10_0: out = 8'b1_11_0_00_11;
        9'b0_11_1_00_10_1: out = 8'b1_11_0_00_11;
        9'b0_11_1_00_11_0: out = 8'b1_10_0_01_11;
        9'b0_11_1_00_11_1: out = 8'b1_01_0_10_11;
        9'b0_11_1_01_00_0: out = 8'bx_xx_x_xx_xx;
        9'b0_11_1_01_00_1: out = 8'bx_xx_x_xx_xx;
        9'b0_11_1_01_01_0: out = 8'bx_xx_x_xx_xx;
        9'b0_11_1_01_01_1: out = 8'bx_xx_x_xx_xx;
        9'b0_11_1_01_10_0: out = 8'bx_xx_x_xx_xx;
        9'b0_11_1_01_10_1: out = 8'bx_xx_x_xx_xx;
        9'b0_11_1_01_11_0: out = 8'bx_xx_x_xx_xx;
        9'b0_11_1_01_11_1: out = 8'bx_xx_x_xx_xx;
        9'b0_11_1_10_00_0: out = 8'bx_xx_x_xx_xx;
        9'b0_11_1_10_00_1: out = 8'bx_xx_x_xx_xx;
        9'b0_11_1_10_01_0: out = 8'bx_xx_x_xx_xx;
        9'b0_11_1_10_01_1: out = 8'bx_xx_x_xx_xx;
        9'b0_11_1_10_10_0: out = 8'bx_xx_x_xx_xx;
        9'b0_11_1_10_10_1: out = 8'bx_xx_x_xx_xx;
        9'b0_11_1_10_11_0: out = 8'bx_xx_x_xx_xx;
        9'b0_11_1_10_11_1: out = 8'bx_xx_x_xx_xx;
        9'b0_11_1_11_00_0: out = 8'bx_xx_x_xx_xx;
        9'b0_11_1_11_00_1: out = 8'bx_xx_x_xx_xx;
        9'b0_11_1_11_01_0: out = 8'bx_xx_x_xx_xx;
        9'b0_11_1_11_01_1: out = 8'bx_xx_x_xx_xx;
        9'b0_11_1_11_10_0: out = 8'bx_xx_x_xx_xx;
        9'b0_11_1_11_10_1: out = 8'bx_xx_x_xx_xx;
        9'b0_11_1_11_11_0: out = 8'bx_xx_x_xx_xx;
        9'b0_11_1_11_11_1: out = 8'bx_xx_x_xx_xx;
        9'b1_00_0_00_00_0: out = 8'b1_00_0_00_00;
        9'b1_00_0_00_00_1: out = 8'b1_00_0_00_00;
        9'b1_00_0_00_01_0: out = 8'b1_00_0_00_00;
        9'b1_00_0_00_01_1: out = 8'b1_00_0_00_00;
        9'b1_00_0_00_10_0: out = 8'b1_00_0_00_00;
        9'b1_00_0_00_10_1: out = 8'b1_00_0_00_00;
        9'b1_00_0_00_11_0: out = 8'b1_00_0_00_00;
        9'b1_00_0_00_11_1: out = 8'b1_00_0_00_00;
        9'b1_00_0_01_00_0: out = 8'b1_01_0_00_01;
        9'b1_00_0_01_00_1: out = 8'b1_00_0_01_01;
        9'b1_00_0_01_01_0: out = 8'b1_00_0_01_00;
        9'b1_00_0_01_01_1: out = 8'b1_00_0_01_00;
        9'b1_00_0_01_10_0: out = 8'b1_00_0_01_00;
        9'b1_00_0_01_10_1: out = 8'b1_00_0_01_00;
        9'b1_00_0_01_11_0: out = 8'b1_00_0_01_00;
        9'b1_00_0_01_11_1: out = 8'b1_00_0_01_00;
        9'b1_00_0_10_00_0: out = 8'b1_10_0_00_01;
        9'b1_00_0_10_00_1: out = 8'b1_01_0_01_01;
        9'b1_00_0_10_01_0: out = 8'b1_00_0_10_00;
        9'b1_00_0_10_01_1: out = 8'b1_00_0_10_00;
        9'b1_00_0_10_10_0: out = 8'b1_00_0_10_00;
        9'b1_00_0_10_10_1: out = 8'b1_00_0_10_00;
        9'b1_00_0_10_11_0: out = 8'b1_00_0_10_00;
        9'b1_00_0_10_11_1: out = 8'b1_00_0_10_00;
        9'b1_00_0_11_00_0: out = 8'b1_10_0_01_01;
        9'b1_00_0_11_00_1: out = 8'b1_01_0_10_01;
        9'b1_00_0_11_01_0: out = 8'b1_00_0_11_00;
        9'b1_00_0_11_01_1: out = 8'b1_00_0_11_00;
        9'b1_00_0_11_10_0: out = 8'b1_00_0_11_00;
        9'b1_00_0_11_10_1: out = 8'b1_00_0_11_00;
        9'b1_00_0_11_11_0: out = 8'b1_00_0_11_00;
        9'b1_00_0_11_11_1: out = 8'b1_00_0_11_00;
        9'b1_00_1_00_00_0: out = 8'b1_00_1_00_00;
        9'b1_00_1_00_00_1: out = 8'b1_00_1_00_00;
        9'b1_00_1_00_01_0: out = 8'b1_00_1_00_00;
        9'b1_00_1_00_01_1: out = 8'b1_00_1_00_00;
        9'b1_00_1_00_10_0: out = 8'b1_00_1_00_00;
        9'b1_00_1_00_10_1: out = 8'b1_00_1_00_00;
        9'b1_00_1_00_11_0: out = 8'b1_00_1_00_00;
        9'b1_00_1_00_11_1: out = 8'b1_00_1_00_00;
        9'b1_00_1_01_00_0: out = 8'b1_00_1_01_00;
        9'b1_00_1_01_00_1: out = 8'b1_00_1_01_00;
        9'b1_00_1_01_01_0: out = 8'b1_00_1_01_00;
        9'b1_00_1_01_01_1: out = 8'b1_00_1_01_00;
        9'b1_00_1_01_10_0: out = 8'b1_00_1_01_00;
        9'b1_00_1_01_10_1: out = 8'b1_00_1_01_00;
        9'b1_00_1_01_11_0: out = 8'b1_01_1_00_01;
        9'b1_00_1_01_11_1: out = 8'b1_00_1_01_01;
        9'b1_00_1_10_00_0: out = 8'b1_00_1_10_00;
        9'b1_00_1_10_00_1: out = 8'b1_00_1_10_00;
        9'b1_00_1_10_01_0: out = 8'b1_00_1_10_00;
        9'b1_00_1_10_01_1: out = 8'b1_00_1_10_00;
        9'b1_00_1_10_10_0: out = 8'b1_00_1_10_00;
        9'b1_00_1_10_10_1: out = 8'b1_00_1_10_00;
        9'b1_00_1_10_11_0: out = 8'b1_10_1_00_01;
        9'b1_00_1_10_11_1: out = 8'b1_01_1_01_01;
        9'b1_00_1_11_00_0: out = 8'b1_00_1_11_00;
        9'b1_00_1_11_00_1: out = 8'b1_00_1_11_00;
        9'b1_00_1_11_01_0: out = 8'b1_00_1_11_00;
        9'b1_00_1_11_01_1: out = 8'b1_00_1_11_00;
        9'b1_00_1_11_10_0: out = 8'b1_00_1_11_00;
        9'b1_00_1_11_10_1: out = 8'b1_00_1_11_00;
        9'b1_00_1_11_11_0: out = 8'b1_10_1_01_01;
        9'b1_00_1_11_11_1: out = 8'b1_01_1_10_01;
        9'b1_01_0_00_00_0: out = 8'b1_01_0_00_00;
        9'b1_01_0_00_00_1: out = 8'b1_00_0_01_00;
        9'b1_01_0_00_01_0: out = 8'b1_01_0_00_00;
        9'b1_01_0_00_01_1: out = 8'b1_00_0_01_00;
        9'b1_01_0_00_10_0: out = 8'b1_01_0_00_00;
        9'b1_01_0_00_10_1: out = 8'b1_00_0_01_00;
        9'b1_01_0_00_11_0: out = 8'b1_01_0_00_00;
        9'b1_01_0_00_11_1: out = 8'b1_00_0_01_00;
        9'b1_01_0_01_00_0: out = 8'b1_01_0_01_00;
        9'b1_01_0_01_00_1: out = 8'b1_00_0_10_00;
        9'b1_01_0_01_01_0: out = 8'b1_01_0_01_00;
        9'b1_01_0_01_01_1: out = 8'b1_00_0_10_00;
        9'b1_01_0_01_10_0: out = 8'b1_01_0_01_00;
        9'b1_01_0_01_10_1: out = 8'b1_00_0_10_00;
        9'b1_01_0_01_11_0: out = 8'b1_01_0_01_00;
        9'b1_01_0_01_11_1: out = 8'b1_00_0_10_00;
        9'b1_01_0_10_00_0: out = 8'b1_01_0_10_00;
        9'b1_01_0_10_00_1: out = 8'b1_00_0_11_00;
        9'b1_01_0_10_01_0: out = 8'b1_01_0_10_00;
        9'b1_01_0_10_01_1: out = 8'b1_00_0_11_00;
        9'b1_01_0_10_10_0: out = 8'b1_01_0_10_00;
        9'b1_01_0_10_10_1: out = 8'b1_00_0_11_00;
        9'b1_01_0_10_11_0: out = 8'b1_01_0_10_00;
        9'b1_01_0_10_11_1: out = 8'b1_00_0_11_00;
        9'b1_01_0_11_00_0: out = 8'bx_xx_x_xx_xx;
        9'b1_01_0_11_00_1: out = 8'bx_xx_x_xx_xx;
        9'b1_01_0_11_01_0: out = 8'bx_xx_x_xx_xx;
        9'b1_01_0_11_01_1: out = 8'bx_xx_x_xx_xx;
        9'b1_01_0_11_10_0: out = 8'bx_xx_x_xx_xx;
        9'b1_01_0_11_10_1: out = 8'bx_xx_x_xx_xx;
        9'b1_01_0_11_11_0: out = 8'bx_xx_x_xx_xx;
        9'b1_01_0_11_11_1: out = 8'bx_xx_x_xx_xx;
        9'b1_01_1_00_00_0: out = 8'b1_01_1_00_00;
        9'b1_01_1_00_00_1: out = 8'b1_00_1_01_00;
        9'b1_01_1_00_01_0: out = 8'b1_01_1_00_00;
        9'b1_01_1_00_01_1: out = 8'b1_00_1_01_00;
        9'b1_01_1_00_10_0: out = 8'b1_01_1_00_00;
        9'b1_01_1_00_10_1: out = 8'b1_00_1_01_00;
        9'b1_01_1_00_11_0: out = 8'b1_01_1_00_00;
        9'b1_01_1_00_11_1: out = 8'b1_00_1_01_00;
        9'b1_01_1_01_00_0: out = 8'b1_01_1_01_00;
        9'b1_01_1_01_00_1: out = 8'b1_00_1_10_00;
        9'b1_01_1_01_01_0: out = 8'b1_01_1_01_00;
        9'b1_01_1_01_01_1: out = 8'b1_00_1_10_00;
        9'b1_01_1_01_10_0: out = 8'b1_01_1_01_00;
        9'b1_01_1_01_10_1: out = 8'b1_00_1_10_00;
        9'b1_01_1_01_11_0: out = 8'b1_01_1_01_00;
        9'b1_01_1_01_11_1: out = 8'b1_00_1_10_00;
        9'b1_01_1_10_00_0: out = 8'b1_01_1_10_00;
        9'b1_01_1_10_00_1: out = 8'b1_00_1_11_00;
        9'b1_01_1_10_01_0: out = 8'b1_01_1_10_00;
        9'b1_01_1_10_01_1: out = 8'b1_00_1_11_00;
        9'b1_01_1_10_10_0: out = 8'b1_01_1_10_00;
        9'b1_01_1_10_10_1: out = 8'b1_00_1_11_00;
        9'b1_01_1_10_11_0: out = 8'b1_01_1_10_00;
        9'b1_01_1_10_11_1: out = 8'b1_00_1_11_00;
        9'b1_01_1_11_00_0: out = 8'bx_xx_x_xx_xx;
        9'b1_01_1_11_00_1: out = 8'bx_xx_x_xx_xx;
        9'b1_01_1_11_01_0: out = 8'bx_xx_x_xx_xx;
        9'b1_01_1_11_01_1: out = 8'bx_xx_x_xx_xx;
        9'b1_01_1_11_10_0: out = 8'bx_xx_x_xx_xx;
        9'b1_01_1_11_10_1: out = 8'bx_xx_x_xx_xx;
        9'b1_01_1_11_11_0: out = 8'bx_xx_x_xx_xx;
        9'b1_01_1_11_11_1: out = 8'bx_xx_x_xx_xx;
        9'b1_10_0_00_00_0: out = 8'b1_10_0_00_00;
        9'b1_10_0_00_00_1: out = 8'b1_10_0_00_00;
        9'b1_10_0_00_01_0: out = 8'b1_10_0_00_00;
        9'b1_10_0_00_01_1: out = 8'b1_10_0_00_00;
        9'b1_10_0_00_10_0: out = 8'b1_10_0_00_00;
        9'b1_10_0_00_10_1: out = 8'b1_10_0_00_00;
        9'b1_10_0_00_11_0: out = 8'b1_10_0_00_00;
        9'b1_10_0_00_11_1: out = 8'b1_10_0_00_00;
        9'b1_10_0_01_00_0: out = 8'b1_11_0_00_00;
        9'b1_10_0_01_00_1: out = 8'b1_10_0_01_00;
        9'b1_10_0_01_01_0: out = 8'b1_11_0_00_00;
        9'b1_10_0_01_01_1: out = 8'b1_10_0_01_00;
        9'b1_10_0_01_10_0: out = 8'b1_11_0_00_00;
        9'b1_10_0_01_10_1: out = 8'b1_10_0_01_00;
        9'b1_10_0_01_11_0: out = 8'b1_11_0_00_00;
        9'b1_10_0_01_11_1: out = 8'b1_10_0_01_00;
        9'b1_10_0_10_00_0: out = 8'bx_xx_x_xx_xx;
        9'b1_10_0_10_00_1: out = 8'bx_xx_x_xx_xx;
        9'b1_10_0_10_01_0: out = 8'bx_xx_x_xx_xx;
        9'b1_10_0_10_01_1: out = 8'bx_xx_x_xx_xx;
        9'b1_10_0_10_10_0: out = 8'bx_xx_x_xx_xx;
        9'b1_10_0_10_10_1: out = 8'bx_xx_x_xx_xx;
        9'b1_10_0_10_11_0: out = 8'bx_xx_x_xx_xx;
        9'b1_10_0_10_11_1: out = 8'bx_xx_x_xx_xx;
        9'b1_10_0_11_00_0: out = 8'bx_xx_x_xx_xx;
        9'b1_10_0_11_00_1: out = 8'bx_xx_x_xx_xx;
        9'b1_10_0_11_01_0: out = 8'bx_xx_x_xx_xx;
        9'b1_10_0_11_01_1: out = 8'bx_xx_x_xx_xx;
        9'b1_10_0_11_10_0: out = 8'bx_xx_x_xx_xx;
        9'b1_10_0_11_10_1: out = 8'bx_xx_x_xx_xx;
        9'b1_10_0_11_11_0: out = 8'bx_xx_x_xx_xx;
        9'b1_10_0_11_11_1: out = 8'bx_xx_x_xx_xx;
        9'b1_10_1_00_00_0: out = 8'b1_10_1_00_00;
        9'b1_10_1_00_00_1: out = 8'b1_10_1_00_00;
        9'b1_10_1_00_01_0: out = 8'b1_10_1_00_00;
        9'b1_10_1_00_01_1: out = 8'b1_10_1_00_00;
        9'b1_10_1_00_10_0: out = 8'b1_10_1_00_00;
        9'b1_10_1_00_10_1: out = 8'b1_10_1_00_00;
        9'b1_10_1_00_11_0: out = 8'b1_10_1_00_00;
        9'b1_10_1_00_11_1: out = 8'b1_10_1_00_00;
        9'b1_10_1_01_00_0: out = 8'b1_11_1_00_00;
        9'b1_10_1_01_00_1: out = 8'b1_10_1_01_00;
        9'b1_10_1_01_01_0: out = 8'b1_11_1_00_00;
        9'b1_10_1_01_01_1: out = 8'b1_10_1_01_00;
        9'b1_10_1_01_10_0: out = 8'b1_11_1_00_00;
        9'b1_10_1_01_10_1: out = 8'b1_10_1_01_00;
        9'b1_10_1_01_11_0: out = 8'b1_11_1_00_00;
        9'b1_10_1_01_11_1: out = 8'b1_10_1_01_00;
        9'b1_10_1_10_00_0: out = 8'bx_xx_x_xx_xx;
        9'b1_10_1_10_00_1: out = 8'bx_xx_x_xx_xx;
        9'b1_10_1_10_01_0: out = 8'bx_xx_x_xx_xx;
        9'b1_10_1_10_01_1: out = 8'bx_xx_x_xx_xx;
        9'b1_10_1_10_10_0: out = 8'bx_xx_x_xx_xx;
        9'b1_10_1_10_10_1: out = 8'bx_xx_x_xx_xx;
        9'b1_10_1_10_11_0: out = 8'bx_xx_x_xx_xx;
        9'b1_10_1_10_11_1: out = 8'bx_xx_x_xx_xx;
        9'b1_10_1_11_00_0: out = 8'bx_xx_x_xx_xx;
        9'b1_10_1_11_00_1: out = 8'bx_xx_x_xx_xx;
        9'b1_10_1_11_01_0: out = 8'bx_xx_x_xx_xx;
        9'b1_10_1_11_01_1: out = 8'bx_xx_x_xx_xx;
        9'b1_10_1_11_10_0: out = 8'bx_xx_x_xx_xx;
        9'b1_10_1_11_10_1: out = 8'bx_xx_x_xx_xx;
        9'b1_10_1_11_11_0: out = 8'bx_xx_x_xx_xx;
        9'b1_10_1_11_11_1: out = 8'bx_xx_x_xx_xx;
        9'b1_11_0_00_00_0: out = 8'b1_11_0_00_00;
        9'b1_11_0_00_00_1: out = 8'b1_11_0_00_00;
        9'b1_11_0_00_01_0: out = 8'b1_11_0_00_00;
        9'b1_11_0_00_01_1: out = 8'b1_11_0_00_00;
        9'b1_11_0_00_10_0: out = 8'b1_11_0_00_00;
        9'b1_11_0_00_10_1: out = 8'b1_11_0_00_00;
        9'b1_11_0_00_11_0: out = 8'b1_11_0_00_00;
        9'b1_11_0_00_11_1: out = 8'b1_11_0_00_00;
        9'b1_11_0_01_00_0: out = 8'bx_xx_x_xx_xx;
        9'b1_11_0_01_00_1: out = 8'bx_xx_x_xx_xx;
        9'b1_11_0_01_01_0: out = 8'bx_xx_x_xx_xx;
        9'b1_11_0_01_01_1: out = 8'bx_xx_x_xx_xx;
        9'b1_11_0_01_10_0: out = 8'bx_xx_x_xx_xx;
        9'b1_11_0_01_10_1: out = 8'bx_xx_x_xx_xx;
        9'b1_11_0_01_11_0: out = 8'bx_xx_x_xx_xx;
        9'b1_11_0_01_11_1: out = 8'bx_xx_x_xx_xx;
        9'b1_11_0_10_00_0: out = 8'bx_xx_x_xx_xx;
        9'b1_11_0_10_00_1: out = 8'bx_xx_x_xx_xx;
        9'b1_11_0_10_01_0: out = 8'bx_xx_x_xx_xx;
        9'b1_11_0_10_01_1: out = 8'bx_xx_x_xx_xx;
        9'b1_11_0_10_10_0: out = 8'bx_xx_x_xx_xx;
        9'b1_11_0_10_10_1: out = 8'bx_xx_x_xx_xx;
        9'b1_11_0_10_11_0: out = 8'bx_xx_x_xx_xx;
        9'b1_11_0_10_11_1: out = 8'bx_xx_x_xx_xx;
        9'b1_11_0_11_00_0: out = 8'bx_xx_x_xx_xx;
        9'b1_11_0_11_00_1: out = 8'bx_xx_x_xx_xx;
        9'b1_11_0_11_01_0: out = 8'bx_xx_x_xx_xx;
        9'b1_11_0_11_01_1: out = 8'bx_xx_x_xx_xx;
        9'b1_11_0_11_10_0: out = 8'bx_xx_x_xx_xx;
        9'b1_11_0_11_10_1: out = 8'bx_xx_x_xx_xx;
        9'b1_11_0_11_11_0: out = 8'bx_xx_x_xx_xx;
        9'b1_11_0_11_11_1: out = 8'bx_xx_x_xx_xx;
        9'b1_11_1_00_00_0: out = 8'b1_11_1_00_00;
        9'b1_11_1_00_00_1: out = 8'b1_11_1_00_00;
        9'b1_11_1_00_01_0: out = 8'b1_11_1_00_00;
        9'b1_11_1_00_01_1: out = 8'b1_11_1_00_00;
        9'b1_11_1_00_10_0: out = 8'b1_11_1_00_00;
        9'b1_11_1_00_10_1: out = 8'b1_11_1_00_00;
        9'b1_11_1_00_11_0: out = 8'b1_11_1_00_00;
        9'b1_11_1_00_11_1: out = 8'b1_11_1_00_00;
        9'b1_11_1_01_00_0: out = 8'bx_xx_x_xx_xx;
        9'b1_11_1_01_00_1: out = 8'bx_xx_x_xx_xx;
        9'b1_11_1_01_01_0: out = 8'bx_xx_x_xx_xx;
        9'b1_11_1_01_01_1: out = 8'bx_xx_x_xx_xx;
        9'b1_11_1_01_10_0: out = 8'bx_xx_x_xx_xx;
        9'b1_11_1_01_10_1: out = 8'bx_xx_x_xx_xx;
        9'b1_11_1_01_11_0: out = 8'bx_xx_x_xx_xx;
        9'b1_11_1_01_11_1: out = 8'bx_xx_x_xx_xx;
        9'b1_11_1_10_00_0: out = 8'bx_xx_x_xx_xx;
        9'b1_11_1_10_00_1: out = 8'bx_xx_x_xx_xx;
        9'b1_11_1_10_01_0: out = 8'bx_xx_x_xx_xx;
        9'b1_11_1_10_01_1: out = 8'bx_xx_x_xx_xx;
        9'b1_11_1_10_10_0: out = 8'bx_xx_x_xx_xx;
        9'b1_11_1_10_10_1: out = 8'bx_xx_x_xx_xx;
        9'b1_11_1_10_11_0: out = 8'bx_xx_x_xx_xx;
        9'b1_11_1_10_11_1: out = 8'bx_xx_x_xx_xx;
        9'b1_11_1_11_00_0: out = 8'bx_xx_x_xx_xx;
        9'b1_11_1_11_00_1: out = 8'bx_xx_x_xx_xx;
        9'b1_11_1_11_01_0: out = 8'bx_xx_x_xx_xx;
        9'b1_11_1_11_01_1: out = 8'bx_xx_x_xx_xx;
        9'b1_11_1_11_10_0: out = 8'bx_xx_x_xx_xx;
        9'b1_11_1_11_10_1: out = 8'bx_xx_x_xx_xx;
        9'b1_11_1_11_11_0: out = 8'bx_xx_x_xx_xx;
        9'b1_11_1_11_11_1: out = 8'bx_xx_x_xx_xx;
    endcase
end

endmodule
