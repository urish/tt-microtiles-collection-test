module logo_table(
		input wire [9:0] addr,
		output wire data
	);

	reg d;
	always @(*) begin
		case (addr)
			0: d = 0;
			1: d = 0;
			2: d = 0;
			3: d = 0;
			4: d = 0;
			5: d = 0;
			6: d = 0;
			7: d = 0;
			8: d = 1;
			9: d = 0;
			10: d = 1;
			11: d = 1;
			12: d = 1;
			13: d = 1;
			14: d = 0;
			15: d = 0;
			16: d = 0;
			17: d = 0;
			18: d = 0;
			19: d = 0;
			20: d = 0;
			21: d = 0;
			22: d = 0;
			23: d = 0;
			24: d = 0;
			25: d = 0;
			26: d = 0;
			27: d = 0;
			28: d = 1;
			29: d = 0;
			30: d = 0;
			31: d = 0;
			32: d = 0;
			33: d = 0;
			34: d = 0;
			35: d = 0;
			36: d = 0;
			37: d = 0;
			38: d = 1;
			39: d = 0;
			40: d = 0;
			41: d = 0;
			42: d = 1;
			43: d = 0;
			44: d = 0;
			45: d = 1;
			46: d = 0;
			47: d = 0;
			48: d = 0;
			49: d = 0;
			50: d = 0;
			51: d = 0;
			52: d = 0;
			53: d = 0;
			54: d = 0;
			55: d = 0;
			56: d = 0;
			57: d = 0;
			58: d = 1;
			59: d = 0;
			60: d = 1;
			61: d = 1;
			62: d = 0;
			63: d = 0;
			64: d = 0;
			65: d = 0;
			66: d = 0;
			67: d = 0;
			68: d = 1;
			69: d = 0;
			70: d = 1;
			71: d = 1;
			72: d = 1;
			73: d = 0;
			74: d = 0;
			75: d = 1;
			76: d = 1;
			77: d = 0;
			78: d = 0;
			79: d = 0;
			80: d = 0;
			81: d = 0;
			82: d = 0;
			83: d = 0;
			84: d = 0;
			85: d = 0;
			86: d = 0;
			87: d = 0;
			88: d = 1;
			89: d = 0;
			90: d = 1;
			91: d = 1;
			92: d = 1;
			93: d = 1;
			94: d = 0;
			95: d = 0;
			96: d = 0;
			97: d = 0;
			98: d = 1;
			99: d = 0;
			100: d = 0;
			101: d = 1;
			102: d = 1;
			103: d = 1;
			104: d = 0;
			105: d = 1;
			106: d = 1;
			107: d = 0;
			108: d = 1;
			109: d = 1;
			110: d = 0;
			111: d = 0;
			112: d = 0;
			113: d = 0;
			114: d = 0;
			115: d = 0;
			116: d = 0;
			117: d = 0;
			118: d = 1;
			119: d = 0;
			120: d = 0;
			121: d = 0;
			122: d = 1;
			123: d = 0;
			124: d = 0;
			125: d = 1;
			126: d = 0;
			127: d = 0;
			128: d = 0;
			129: d = 0;
			130: d = 1;
			131: d = 1;
			132: d = 0;
			133: d = 0;
			134: d = 0;
			135: d = 0;
			136: d = 1;
			137: d = 0;
			138: d = 0;
			139: d = 1;
			140: d = 0;
			141: d = 1;
			142: d = 0;
			143: d = 0;
			144: d = 0;
			145: d = 0;
			146: d = 0;
			147: d = 0;
			148: d = 1;
			149: d = 0;
			150: d = 1;
			151: d = 1;
			152: d = 1;
			153: d = 0;
			154: d = 0;
			155: d = 1;
			156: d = 1;
			157: d = 0;
			158: d = 0;
			159: d = 0;
			160: d = 0;
			161: d = 0;
			162: d = 1;
			163: d = 1;
			164: d = 0;
			165: d = 1;
			166: d = 1;
			167: d = 0;
			168: d = 1;
			169: d = 1;
			170: d = 0;
			171: d = 0;
			172: d = 0;
			173: d = 0;
			174: d = 0;
			175: d = 0;
			176: d = 0;
			177: d = 0;
			178: d = 1;
			179: d = 0;
			180: d = 0;
			181: d = 1;
			182: d = 1;
			183: d = 1;
			184: d = 0;
			185: d = 1;
			186: d = 1;
			187: d = 0;
			188: d = 0;
			189: d = 1;
			190: d = 0;
			191: d = 0;
			192: d = 0;
			193: d = 0;
			194: d = 0;
			195: d = 1;
			196: d = 1;
			197: d = 0;
			198: d = 0;
			199: d = 1;
			200: d = 0;
			201: d = 1;
			202: d = 1;
			203: d = 0;
			204: d = 1;
			205: d = 1;
			206: d = 0;
			207: d = 0;
			208: d = 0;
			209: d = 0;
			210: d = 1;
			211: d = 1;
			212: d = 0;
			213: d = 0;
			214: d = 0;
			215: d = 0;
			216: d = 1;
			217: d = 0;
			218: d = 0;
			219: d = 1;
			220: d = 1;
			221: d = 0;
			222: d = 0;
			223: d = 0;
			224: d = 0;
			225: d = 0;
			226: d = 0;
			227: d = 0;
			228: d = 1;
			229: d = 1;
			230: d = 0;
			231: d = 0;
			232: d = 1;
			233: d = 0;
			234: d = 0;
			235: d = 1;
			236: d = 1;
			237: d = 1;
			238: d = 0;
			239: d = 0;
			240: d = 0;
			241: d = 0;
			242: d = 1;
			243: d = 1;
			244: d = 0;
			245: d = 1;
			246: d = 1;
			247: d = 0;
			248: d = 1;
			249: d = 1;
			250: d = 1;
			251: d = 0;
			252: d = 0;
			253: d = 1;
			254: d = 0;
			255: d = 0;
			256: d = 0;
			257: d = 0;
			258: d = 0;
			259: d = 0;
			260: d = 0;
			261: d = 1;
			262: d = 1;
			263: d = 0;
			264: d = 0;
			265: d = 1;
			266: d = 1;
			267: d = 1;
			268: d = 1;
			269: d = 1;
			270: d = 0;
			271: d = 0;
			272: d = 0;
			273: d = 0;
			274: d = 0;
			275: d = 1;
			276: d = 1;
			277: d = 0;
			278: d = 0;
			279: d = 1;
			280: d = 1;
			281: d = 1;
			282: d = 0;
			283: d = 1;
			284: d = 1;
			285: d = 0;
			286: d = 0;
			287: d = 0;
			288: d = 0;
			289: d = 0;
			290: d = 0;
			291: d = 0;
			292: d = 1;
			293: d = 0;
			294: d = 0;
			295: d = 1;
			296: d = 1;
			297: d = 0;
			298: d = 0;
			299: d = 1;
			300: d = 0;
			301: d = 0;
			302: d = 0;
			303: d = 0;
			304: d = 0;
			305: d = 0;
			306: d = 0;
			307: d = 0;
			308: d = 0;
			309: d = 1;
			310: d = 1;
			311: d = 0;
			312: d = 0;
			313: d = 1;
			314: d = 1;
			315: d = 0;
			316: d = 0;
			317: d = 1;
			318: d = 0;
			319: d = 0;
			320: d = 0;
			321: d = 0;
			322: d = 0;
			323: d = 0;
			324: d = 1;
			325: d = 1;
			326: d = 1;
			327: d = 1;
			328: d = 0;
			329: d = 1;
			330: d = 1;
			331: d = 0;
			332: d = 1;
			333: d = 1;
			334: d = 0;
			335: d = 0;
			336: d = 0;
			337: d = 0;
			338: d = 0;
			339: d = 0;
			340: d = 1;
			341: d = 0;
			342: d = 0;
			343: d = 1;
			344: d = 1;
			345: d = 0;
			346: d = 1;
			347: d = 1;
			348: d = 1;
			349: d = 1;
			350: d = 0;
			351: d = 0;
			352: d = 0;
			353: d = 0;
			354: d = 0;
			355: d = 0;
			356: d = 1;
			357: d = 1;
			358: d = 0;
			359: d = 1;
			360: d = 1;
			361: d = 0;
			362: d = 0;
			363: d = 1;
			364: d = 1;
			365: d = 1;
			366: d = 0;
			367: d = 0;
			368: d = 0;
			369: d = 0;
			370: d = 0;
			371: d = 0;
			372: d = 0;
			373: d = 1;
			374: d = 0;
			375: d = 0;
			376: d = 0;
			377: d = 0;
			378: d = 0;
			379: d = 0;
			380: d = 0;
			381: d = 0;
			382: d = 0;
			383: d = 0;
			384: d = 0;
			385: d = 0;
			386: d = 0;
			387: d = 0;
			388: d = 0;
			389: d = 0;
			390: d = 1;
			391: d = 0;
			392: d = 0;
			393: d = 1;
			394: d = 1;
			395: d = 0;
			396: d = 0;
			397: d = 1;
			398: d = 0;
			399: d = 0;
			400: d = 0;
			401: d = 0;
			402: d = 0;
			403: d = 0;
			404: d = 1;
			405: d = 0;
			406: d = 1;
			407: d = 1;
			408: d = 1;
			409: d = 1;
			410: d = 1;
			411: d = 1;
			412: d = 0;
			413: d = 1;
			414: d = 0;
			415: d = 0;
			416: d = 0;
			417: d = 0;
			418: d = 0;
			419: d = 0;
			420: d = 1;
			421: d = 0;
			422: d = 0;
			423: d = 1;
			424: d = 1;
			425: d = 0;
			426: d = 0;
			427: d = 1;
			428: d = 1;
			429: d = 0;
			430: d = 0;
			431: d = 0;
			432: d = 0;
			433: d = 0;
			434: d = 0;
			435: d = 0;
			436: d = 1;
			437: d = 1;
			438: d = 0;
			439: d = 0;
			440: d = 1;
			441: d = 0;
			442: d = 0;
			443: d = 1;
			444: d = 0;
			445: d = 0;
			446: d = 0;
			447: d = 0;
			448: d = 0;
			449: d = 0;
			450: d = 0;
			451: d = 0;
			452: d = 0;
			453: d = 1;
			454: d = 1;
			455: d = 0;
			456: d = 0;
			457: d = 1;
			458: d = 1;
			459: d = 0;
			460: d = 1;
			461: d = 1;
			462: d = 0;
			463: d = 0;
			464: d = 0;
			465: d = 0;
			466: d = 0;
			467: d = 0;
			468: d = 1;
			469: d = 1;
			470: d = 1;
			471: d = 1;
			472: d = 0;
			473: d = 1;
			474: d = 1;
			475: d = 0;
			476: d = 1;
			477: d = 1;
			478: d = 0;
			479: d = 0;
			480: d = 0;
			481: d = 0;
			482: d = 0;
			483: d = 0;
			484: d = 1;
			485: d = 0;
			486: d = 0;
			487: d = 1;
			488: d = 1;
			489: d = 0;
			490: d = 0;
			491: d = 1;
			492: d = 0;
			493: d = 1;
			494: d = 0;
			495: d = 0;
			496: d = 0;
			497: d = 0;
			498: d = 0;
			499: d = 0;
			500: d = 1;
			501: d = 1;
			502: d = 0;
			503: d = 1;
			504: d = 1;
			505: d = 0;
			506: d = 0;
			507: d = 1;
			508: d = 1;
			509: d = 1;
			510: d = 0;
			511: d = 0;
			512: d = 0;
			513: d = 0;
			514: d = 0;
			515: d = 0;
			516: d = 0;
			517: d = 1;
			518: d = 1;
			519: d = 0;
			520: d = 1;
			521: d = 1;
			522: d = 0;
			523: d = 0;
			524: d = 1;
			525: d = 0;
			526: d = 0;
			527: d = 0;
			528: d = 0;
			529: d = 0;
			530: d = 0;
			531: d = 0;
			532: d = 0;
			533: d = 0;
			534: d = 1;
			535: d = 0;
			536: d = 0;
			537: d = 1;
			538: d = 1;
			539: d = 0;
			540: d = 0;
			541: d = 1;
			542: d = 0;
			543: d = 0;
			544: d = 0;
			545: d = 0;
			546: d = 0;
			547: d = 0;
			548: d = 1;
			549: d = 0;
			550: d = 0;
			551: d = 1;
			552: d = 0;
			553: d = 1;
			554: d = 1;
			555: d = 0;
			556: d = 0;
			557: d = 1;
			558: d = 0;
			559: d = 0;
			560: d = 0;
			561: d = 0;
			562: d = 0;
			563: d = 0;
			564: d = 1;
			565: d = 0;
			566: d = 0;
			567: d = 1;
			568: d = 1;
			569: d = 0;
			570: d = 0;
			571: d = 1;
			572: d = 0;
			573: d = 0;
			574: d = 0;
			575: d = 0;
			576: d = 0;
			577: d = 0;
			578: d = 0;
			579: d = 0;
			580: d = 1;
			581: d = 1;
			582: d = 0;
			583: d = 0;
			584: d = 1;
			585: d = 0;
			586: d = 0;
			587: d = 1;
			588: d = 0;
			589: d = 0;
			590: d = 0;
			591: d = 0;
			592: d = 0;
			593: d = 0;
			594: d = 0;
			595: d = 0;
			596: d = 1;
			597: d = 1;
			598: d = 1;
			599: d = 1;
			600: d = 0;
			601: d = 1;
			602: d = 1;
			603: d = 0;
			604: d = 1;
			605: d = 1;
			606: d = 0;
			607: d = 0;
			608: d = 0;
			609: d = 0;
			610: d = 0;
			611: d = 0;
			612: d = 1;
			613: d = 1;
			614: d = 1;
			615: d = 0;
			616: d = 1;
			617: d = 1;
			618: d = 1;
			619: d = 1;
			620: d = 0;
			621: d = 1;
			622: d = 0;
			623: d = 0;
			624: d = 0;
			625: d = 0;
			626: d = 0;
			627: d = 0;
			628: d = 1;
			629: d = 1;
			630: d = 0;
			631: d = 1;
			632: d = 1;
			633: d = 0;
			634: d = 0;
			635: d = 1;
			636: d = 1;
			637: d = 1;
			638: d = 0;
			639: d = 0;
			640: d = 0;
			641: d = 0;
			642: d = 0;
			643: d = 0;
			644: d = 0;
			645: d = 1;
			646: d = 0;
			647: d = 0;
			648: d = 1;
			649: d = 0;
			650: d = 0;
			651: d = 1;
			652: d = 1;
			653: d = 0;
			654: d = 0;
			655: d = 0;
			656: d = 0;
			657: d = 0;
			658: d = 0;
			659: d = 0;
			660: d = 0;
			661: d = 0;
			662: d = 1;
			663: d = 0;
			664: d = 0;
			665: d = 1;
			666: d = 1;
			667: d = 0;
			668: d = 1;
			669: d = 1;
			670: d = 0;
			671: d = 0;
			672: d = 0;
			673: d = 0;
			674: d = 0;
			675: d = 0;
			676: d = 1;
			677: d = 0;
			678: d = 1;
			679: d = 0;
			680: d = 0;
			681: d = 1;
			682: d = 1;
			683: d = 0;
			684: d = 0;
			685: d = 1;
			686: d = 0;
			687: d = 0;
			688: d = 0;
			689: d = 0;
			690: d = 0;
			691: d = 0;
			692: d = 1;
			693: d = 0;
			694: d = 0;
			695: d = 1;
			696: d = 1;
			697: d = 0;
			698: d = 0;
			699: d = 1;
			700: d = 1;
			701: d = 1;
			702: d = 0;
			703: d = 0;
			704: d = 0;
			705: d = 0;
			706: d = 0;
			707: d = 0;
			708: d = 1;
			709: d = 1;
			710: d = 0;
			711: d = 0;
			712: d = 1;
			713: d = 0;
			714: d = 0;
			715: d = 1;
			716: d = 1;
			717: d = 0;
			718: d = 0;
			719: d = 0;
			720: d = 0;
			721: d = 0;
			722: d = 0;
			723: d = 0;
			724: d = 0;
			725: d = 1;
			726: d = 1;
			727: d = 0;
			728: d = 0;
			729: d = 1;
			730: d = 1;
			731: d = 0;
			732: d = 0;
			733: d = 1;
			734: d = 1;
			735: d = 0;
			736: d = 0;
			737: d = 0;
			738: d = 0;
			739: d = 0;
			740: d = 1;
			741: d = 1;
			742: d = 1;
			743: d = 0;
			744: d = 0;
			745: d = 1;
			746: d = 1;
			747: d = 0;
			748: d = 0;
			749: d = 1;
			750: d = 0;
			751: d = 0;
			752: d = 0;
			753: d = 0;
			754: d = 0;
			755: d = 0;
			756: d = 1;
			757: d = 0;
			758: d = 0;
			759: d = 1;
			760: d = 1;
			761: d = 0;
			762: d = 0;
			763: d = 1;
			764: d = 1;
			765: d = 0;
			766: d = 1;
			767: d = 1;
			768: d = 0;
			769: d = 0;
			770: d = 0;
			771: d = 0;
			772: d = 1;
			773: d = 1;
			774: d = 0;
			775: d = 1;
			776: d = 1;
			777: d = 0;
			778: d = 0;
			779: d = 1;
			780: d = 1;
			781: d = 0;
			782: d = 0;
			783: d = 0;
			784: d = 0;
			785: d = 0;
			786: d = 0;
			787: d = 0;
			788: d = 0;
			789: d = 1;
			790: d = 1;
			791: d = 0;
			792: d = 0;
			793: d = 1;
			794: d = 1;
			795: d = 0;
			796: d = 1;
			797: d = 1;
			798: d = 1;
			799: d = 1;
			800: d = 0;
			801: d = 0;
			802: d = 0;
			803: d = 0;
			804: d = 1;
			805: d = 1;
			806: d = 1;
			807: d = 0;
			808: d = 0;
			809: d = 1;
			810: d = 1;
			811: d = 0;
			812: d = 0;
			813: d = 1;
			814: d = 0;
			815: d = 0;
			816: d = 0;
			817: d = 0;
			818: d = 0;
			819: d = 0;
			820: d = 1;
			821: d = 0;
			822: d = 0;
			823: d = 1;
			824: d = 1;
			825: d = 0;
			826: d = 0;
			827: d = 0;
			828: d = 1;
			829: d = 0;
			830: d = 0;
			831: d = 1;
			832: d = 0;
			833: d = 0;
			834: d = 0;
			835: d = 0;
			836: d = 1;
			837: d = 1;
			838: d = 0;
			839: d = 0;
			840: d = 1;
			841: d = 0;
			842: d = 1;
			843: d = 1;
			844: d = 1;
			845: d = 1;
			846: d = 0;
			847: d = 0;
			848: d = 0;
			849: d = 0;
			850: d = 0;
			851: d = 0;
			852: d = 0;
			853: d = 1;
			854: d = 1;
			855: d = 0;
			856: d = 1;
			857: d = 1;
			858: d = 1;
			859: d = 0;
			860: d = 0;
			861: d = 1;
			862: d = 0;
			863: d = 0;
			864: d = 0;
			865: d = 0;
			866: d = 0;
			867: d = 0;
			868: d = 0;
			869: d = 1;
			870: d = 0;
			871: d = 0;
			872: d = 0;
			873: d = 0;
			874: d = 0;
			875: d = 0;
			876: d = 0;
			877: d = 0;
			878: d = 0;
			879: d = 0;
			880: d = 0;
			881: d = 0;
			882: d = 0;
			883: d = 0;
			884: d = 1;
			885: d = 0;
			886: d = 0;
			887: d = 1;
			888: d = 1;
			889: d = 1;
			890: d = 0;
			891: d = 1;
			892: d = 0;
			893: d = 0;
			894: d = 0;
			895: d = 0;
			896: d = 0;
			897: d = 0;
			898: d = 0;
			899: d = 0;
			900: d = 1;
			901: d = 0;
			902: d = 1;
			903: d = 1;
			904: d = 1;
			905: d = 1;
			906: d = 1;
			907: d = 1;
			908: d = 1;
			909: d = 1;
			910: d = 0;
			911: d = 0;
			912: d = 0;
			913: d = 0;
			914: d = 0;
			915: d = 0;
			916: d = 1;
			917: d = 1;
			918: d = 0;
			919: d = 0;
			920: d = 0;
			921: d = 0;
			922: d = 0;
			923: d = 0;
			924: d = 0;
			925: d = 0;
			926: d = 0;
			927: d = 0;
			928: d = 0;
			929: d = 0;
			930: d = 0;
			931: d = 0;
			932: d = 0;
			933: d = 1;
			934: d = 0;
			935: d = 0;
			936: d = 0;
			937: d = 0;
			938: d = 0;
			939: d = 0;
			940: d = 1;
			941: d = 1;
			942: d = 0;
			943: d = 0;
			944: d = 0;
			945: d = 0;
			946: d = 0;
			947: d = 0;
			948: d = 1;
			949: d = 1;
			950: d = 0;
			951: d = 1;
			952: d = 0;
			953: d = 0;
			954: d = 0;
			955: d = 0;
			956: d = 0;
			957: d = 0;
			958: d = 0;
			959: d = 0;
			960: d = 1'bX;
			961: d = 1'bX;
			962: d = 1'bX;
			963: d = 1'bX;
			964: d = 1'bX;
			965: d = 1'bX;
			966: d = 1'bX;
			967: d = 1'bX;
			968: d = 1'bX;
			969: d = 1'bX;
			970: d = 1'bX;
			971: d = 1'bX;
			972: d = 1'bX;
			973: d = 1'bX;
			974: d = 1'bX;
			975: d = 1'bX;
			976: d = 1'bX;
			977: d = 1'bX;
			978: d = 1'bX;
			979: d = 1'bX;
			980: d = 1'bX;
			981: d = 1'bX;
			982: d = 1'bX;
			983: d = 1'bX;
			984: d = 1'bX;
			985: d = 1'bX;
			986: d = 1'bX;
			987: d = 1'bX;
			988: d = 1'bX;
			989: d = 1'bX;
			990: d = 1'bX;
			991: d = 1'bX;
			992: d = 1'bX;
			993: d = 1'bX;
			994: d = 1'bX;
			995: d = 1'bX;
			996: d = 1'bX;
			997: d = 1'bX;
			998: d = 1'bX;
			999: d = 1'bX;
			1000: d = 1'bX;
			1001: d = 1'bX;
			1002: d = 1'bX;
			1003: d = 1'bX;
			1004: d = 1'bX;
			1005: d = 1'bX;
			1006: d = 1'bX;
			1007: d = 1'bX;
			1008: d = 1'bX;
			1009: d = 1'bX;
			1010: d = 1'bX;
			1011: d = 1'bX;
			1012: d = 1'bX;
			1013: d = 1'bX;
			1014: d = 1'bX;
			1015: d = 1'bX;
			1016: d = 1'bX;
			1017: d = 1'bX;
			1018: d = 1'bX;
			1019: d = 1'bX;
			1020: d = 1'bX;
			1021: d = 1'bX;
			1022: d = 1'bX;
			1023: d = 1'bX;
			default: d = 'X;
		endcase
	end

	assign data = d;
endmodule : logo_table
