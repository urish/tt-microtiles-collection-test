`default_nettype none

module sine_table(
    input wire [4:0] in,
    output reg [11:0] out
);

always @(*) begin
    case(in)
        5'b00000: out = 12'b000001_111111;
        5'b00001: out = 12'b000010_111111;
        5'b00010: out = 12'b000100_111111;
        5'b00011: out = 12'b000101_111111;
        5'b00100: out = 12'b000111_111111;
        5'b00101: out = 12'b001001_111111;
        5'b00110: out = 12'b001010_111111;
        5'b00111: out = 12'b001100_111110;
        5'b01000: out = 12'b001101_111110;
        5'b01001: out = 12'b001111_111110;
        5'b01010: out = 12'b010000_111101;
        5'b01011: out = 12'b010010_111101;
        5'b01100: out = 12'b010011_111101;
        5'b01101: out = 12'b010101_111100;
        5'b01110: out = 12'b010110_111100;
        5'b01111: out = 12'b011000_111011;
        5'b10000: out = 12'b011001_111010;
        5'b10001: out = 12'b011010_111010;
        5'b10010: out = 12'b011100_111001;
        5'b10011: out = 12'b011101_111000;
        5'b10100: out = 12'b011111_111000;
        5'b10101: out = 12'b100000_110111;
        5'b10110: out = 12'b100001_110110;
        5'b10111: out = 12'b100011_110101;
        5'b11000: out = 12'b100100_110100;
        5'b11001: out = 12'b100101_110011;
        5'b11010: out = 12'b100110_110011;
        5'b11011: out = 12'b101000_110010;
        5'b11100: out = 12'b101001_110001;
        5'b11101: out = 12'b101010_110000;
        5'b11110: out = 12'b101011_101111;
        5'b11111: out = 12'b101100_101101;
    endcase
end

endmodule
