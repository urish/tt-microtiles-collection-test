/*
   Verilog module for the inverse AES S-box.

   Copyright 2024 Dag Arne Osvik

   Licensed under the Apache License, Version 2.0 (the "License");
   you may not use this file except in compliance with the License.
   You may obtain a copy of the License at

       http://www.apache.org/licenses/LICENSE-2.0

   Unless required by applicable law or agreed to in writing, software
   distributed under the License is distributed on an "AS IS" BASIS,
   WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
   See the License for the specific language governing permissions and
   limitations under the License.
*/

module sbox_aesinv (
    input            clk,
    input      [7:0] x,
    output     [7:0] y,
    output reg [7:0] cy);

    wire  x55555555;
    wire  x33333333;
    wire  x0f0f0f0f;
    wire  x00ff00ff;
    wire  x0000ffff;

    wire x55;
    wire x33;
    wire x0f;

    assign x55555555 = x[0];
    assign x33333333 = x[1];
    assign x0f0f0f0f = x[2];
    assign x00ff00ff = x[3];
    assign x0000ffff = x[4];

    assign x55 = x[5];
    assign x33 = x[6];
    assign x0f = x[7];

    wire x01;
    wire x02;
    wire x04;
    wire x08;
    wire x10;
    wire x20;
    wire x40;
    wire x80;

    and3 	m01 (.y(x01), .a  (x55), .b  (x33), .c  (x0f));
    and3b 	m02 (.y(x02), .an (x55), .b  (x33), .c  (x0f));
    and3b 	m04 (.y(x04), .an (x33), .b  (x55), .c  (x0f));
    nor3b 	m08 (.y(x08), .an (x0f), .b  (x55), .c  (x33));
    and3b 	m10 (.y(x10), .an (x0f), .b  (x55), .c  (x33));
    nor3b 	m20 (.y(x20), .an (x33), .b  (x55), .c  (x0f));
    nor3b 	m40 (.y(x40), .an (x55), .b  (x33), .c  (x0f));
    nor3 	m80 (.y(x80), .a  (x55), .b  (x33), .c  (x0f));

    wire
        x7, x7a, x7b, x7c, x7d,
        x6, x6a, x6b, x6c, x6d,
        x5, x5a, x5b, x5c, x5d,
        x4, x4a, x4b, x4c, x4d,
        x3, x3a, x3b, x3c, x3d,
        x2, x2a, x2b, x2c, x2d,
        x1, x1a, x1b, x1c, x1d,
        x0, x0a, x0b, x0c, x0d;

    wire x00000008;
    wire x00000013;
    wire x00000054;
    wire x00000080;
    wire x00000117;
    wire x00000550;
    wire x00001011;
    wire x0000101a;
    wire x000010dc;
    wire x00001110;
    wire x00001175;
    wire x00001355;
    wire x00008000;
    wire x00008880;
    wire x0000a000;
    wire x00010005;
    wire x00010031;
    wire x00050011;
    wire x00050022;
    wire x00050300;
    wire x00060006;
    wire x00070013;
    wire x0007173f;
    wire x000a022a;
    wire x000a0808;
    wire x000aaaab;
    wire x000c0e5e;
    wire x000ccc00;
    wire x000f023f;
    wire x00113035;
    wire x00130f0f;
    wire x00330404;
    wire x004000c0;
    wire x005dccdd;
    wire x007fabff;
    wire x0100011f;
    wire x01010003;
    wire x01011010;
    wire x01155fff;
    wire x0133273f;
    wire x0137133f;
    wire x01f731f7;
    wire x03fc03fc;
    wire x04044447;
    wire x040c0000;
    wire x05500000;
    wire x055f0557;
    wire x08000000;
    wire x0a000000;
    wire x0a080000;
    wire x0abf1bbf;
    wire x0b1fafbf;
    wire x0cd37660;
    wire x0e0a0000;
    wire x0eb6ef2f;
    wire x0f5f0a5f;
    wire x0ff7ffff;
    wire x10104040;
    wire x11004400;
    wire x11131313;
    wire x11771333;
    wire x11aa0000;
    wire x12bf5b4f;
    wire x131317df;
    wire x1333131f;
    wire x135f5fdf;
    wire x13bfbfbf;
    wire x15000400;
    wire x151d777f;
    wire x15555050;
    wire x169287dc;
    wire x175f333f;
    wire x17ff555f;
    wire x1a10b72b;
    wire x1d7f5dff;
    wire x1f7b28d7;
    wire x1f7f55ff;
    wire x229616fd;
    wire x23369e29;
    wire x23853f57;
    wire x24cc4461;
    wire x2a000000;
    wire x2aeeaaee;
    wire x2bffafff;
    wire x2c6cdf10;
    wire x2ca62526;
    wire x2d9fb2de;
    wire x2fa5e682;
    wire x2fafffff;
    wire x30307000;
    wire x3030f1f0;
    wire x30c030c0;
    wire x318ab4e1;
    wire x32220000;
    wire x32302020;
    wire x323233fb;
    wire x326fc4dd;
    wire x333300cf;
    wire x33cfffff;
    wire x33ffff0f;
    wire x37303733;
    wire x3777053f;
    wire x37ff5577;
    wire x39fe8cff;
    wire x3c3ffdff;
    wire x3cf25843;
    wire x3f00ff05;
    wire x3f0fffcf;
    wire x3f557fff;
    wire x3fff2faf;
    wire x3fffffff;
    wire x40484048;
    wire x40c00000;
    wire x41d5cc5c;
    wire x4213e265;
    wire x42e28881;
    wire x4332245f;
    wire x434a8cf5;
    wire x43fecdd2;
    wire x4638af86;
    wire x4e5feeff;
    wire x50004000;
    wire x52af6f23;
    wire x52c516d9;
    wire x54eaa319;
    wire x55556666;
    wire x55775071;
    wire x557f00ff;
    wire x571fff3f;
    wire x57ffff00;
    wire x5a5f5b5f;
    wire x5aaa5aaa;
    wire x5b847ba9;
    wire x5e9f51e4;
    wire x5f5ffafa;
    wire x5fff0faf;
    wire x6191ae47;
    wire x6a86145f;
    wire x6ad30f0f;
    wire x6d287e63;
    wire x7077f7ff;
    wire x777717ff;
    wire x77cd77ff;
    wire x77fc77fc;
    wire x77ff3337;
    wire x7847e6db;
    wire x7c7c7c7d;
    wire x7ca10f66;
    wire x7f5f3300;
    wire x80000000;
    wire x80808080;
    wire x854f7ef5;
    wire x88000000;
    wire x88008800;
    wire x88880000;
    wire x88888888;
    wire x8ad2e815;
    wire x8b30445b;
    wire x8df398a3;
    wire x8fdfffff;
    wire x96492239;
    wire x9d97aa84;
    wire xa0008000;
    wire xa000a000;
    wire xa0a00000;
    wire xa0a0a0a0;
    wire xa0a0a1a1;
    wire xa0fb7cd2;
    wire xa1b3a5bf;
    wire xa4b75f65;
    wire xa8000000;
    wire xa8008000;
    wire xa8800000;
    wire xa8a8a8a8;
    wire xa90301b8;
    wire xa9e15289;
    wire xaa000000;
    wire xaa0faf5f;
    wire xaa88aa88;
    wire xaaa0aaa0;
    wire xaaaa0000;
    wire xaaaa8888;
    wire xaaaaa0a0;
    wire xaaaaaa00;
    wire xaaaf153f;
    wire xadffadff;
    wire xaf7faf7f;
    wire xafa5ffff;
    wire xb047c23f;
    wire xb1b1f5f7;
    wire xbb3333ff;
    wire xbb77ffff;
    wire xbbbbf5f5;
    wire xbfbf373f;
    wire xbfffffff;
    wire xc0008000;
    wire xc000c000;
    wire xc011c011;
    wire xc0c00000;
    wire xc0c0c0c0;
    wire xc3c3c3cf;
    wire xc4cf14da;
    wire xc5cfc5df;
    wire xc60b25d3;
    wire xc6aca424;
    wire xc800c000;
    wire xc8c8c8c8;
    wire xcbea0a80;
    wire xcbffcbff;
    wire xcc000000;
    wire xcc00cc00;
    wire xcc880000;
    wire xcc88cc88;
    wire xccc0ccc0;
    wire xcccc0000;
    wire xcccc8888;
    wire xccccc0c0;
    wire xcccccc00;
    wire xcccf030f;
    wire xd1f16c3a;
    wire xd2a0de7f;
    wire xd7997ddd;
    wire xdd11cc00;
    wire xdd5555ff;
    wire xdd7fff7f;
    wire xddf7ddf7;
    wire xdf77df77;
    wire xdfc11244;
    wire xdfdf77ff;
    wire xe080c000;
    wire xe0e0e0e0;
    wire xe2cda26e;
    wire xe3ab5bd2;
    wire xe8133bb7;
    wire xe8e8e800;
    wire xeaeaeaea;
    wire xeaefffff;
    wire xee00ee00;
    wire xeeaaeeaa;
    wire xeecc98e2;
    wire xeeee0000;
    wire xeeee8080;
    wire xeeeeaaaa;
    wire xeeeeeeee;
    wire xef715dd5;
    wire xefefcf8f;
    wire xf0000000;
    wire xf000f000;
    wire xf003f003;
    wire xf0a0a0a0;
    wire xf0a0f0a0;
    wire xf0a0f3a3;
    wire xf0c0c000;
    wire xf0c0f0c0;
    wire xf0c0f5d5;
    wire xf0f00000;
    wire xf0f0a0a0;
    wire xf0f0c0c0;
    wire xf0f0f000;
    wire xf0f0f0f0;
    wire xf12405c2;
    wire xf1a1f1a1;
    wire xf1f1ffff;
    wire xf1f5f5f7;
    wire xf333f377;
    wire xf33fffff;
    wire xf35ff3ff;
    wire xf3f37f7f;
    wire xf446ce08;
    wire xf4bcfdb0;
    wire xf555f57f;
    wire xf5a5ffff;
    wire xf5ff5fff;
    wire xf8008000;
    wire xf8f0c800;
    wire xf8f8c8c8;
    wire xfa00fa00;
    wire xfaaafaaa;
    wire xfac8a080;
    wire xfaf8fa00;
    wire xfafa0000;
    wire xfafaaaaa;
    wire xfafafafa;
    wire xfc00fc00;
    wire xfccca000;
    wire xfcccfccc;
    wire xfccfffff;
    wire xfcecf8a0;
    wire xfcfc0000;
    wire xfcfccccc;
    wire xfcfcccff;
    wire xfcfcf8a0;
    wire xfcfcfcfc;
    wire xfd11ffff;
    wire xfec8eec8;
    wire xfecccc00;
    wire xfeccfec8;
    wire xfeecfaa8;
    wire xfeeef8a8;
    wire xfefaeca8;
    wire xfefafefa;
    wire xfefea8a0;
    wire xfefefefe;
    wire xff000000;
    wire xff00aa00;
    wire xff00cc00;
    wire xff00f000;
    wire xff00ff00;
    wire xff010103;
    wire xff05333f;
    wire xff3f05ff;
    wire xff7f7f7f;
    wire xffaa0000;
    wire xffaaaaaa;
    wire xffaaffaa;
    wire xffb3ffb3;
    wire xffcc0000;
    wire xffcccccc;
    wire xffcceec8;
    wire xffccffcc;
    wire xffddddff;
    wire xffec8888;
    wire xffecece8;
    wire xffecffa8;
    wire xffeeee88;
    wire xffeeffee;
    wire xfff00000;
    wire xfff0f0f0;
    wire xfff0fff0;
    wire xfff30000;
    wire xfff5f5ff;
    wire xfff8fac8;
    wire xfff8ffa0;
    wire xfffafffa;
    wire xfffcfeec;
    wire xfffcfffc;
    wire xfffcfffd;
    wire xfffef888;
    wire xffff0000;
    wire xffff8f0f;
    wire xffffaaaa;
    wire xffffcccc;
    wire xffffeeee;
    wire xfffff0f0;
    wire xfffff8a0;
    wire xfffffafa;
    wire xfffffcfc;
    wire xfffffeee;
    wire xffffff00;
    wire xffffffaa;
    wire xffffffcc;
    wire xffffffdd;
    wire xffffffea;
    wire xffffffec;
    wire xfffffff0;
    wire xfffffffc;
    wire xfffffffe;

    nor2b 	m00000008 (.y(x00000008), .an (xcc88cc88), .b  (xfffffff0));
    nor2 	m00000013 (.y(x00000013), .a  (xf0f0a0a0), .b  (xffffffcc));
    nor2b 	m00000054 (.y(x00000054), .an (xfffffcfc), .b  (xffffffaa));
    nor2b 	m00000080 (.y(x00000080), .an (x80808080), .b  (xf0f0f000));
    nor4 	m00000117 (.y(x00000117), .a  (xffff0000), .b  (xfc00fc00), .c  (xc8c8c8c8), .d  (xaaa0aaa0));
    o22ai 	m00000550 (.y(x00000550), .a0 (x00ff00ff), .a1 (xfffffafa), .b0 (x0f0f0f0f), .b1 (xffffffaa));
    a21oi 	m00001011 (.y(x00001011), .a0 (xff00ff00), .a1 (x0f0f0f0f), .b0 (xffffeeee));
    o22ai 	m0000101a (.y(x0000101a), .a0 (x0f0f0f0f), .a1 (xffffeeee), .b0 (x55555555), .b1 (xfffffff0));
    o22ai 	m000010dc (.y(x000010dc), .a0 (x0f0f0f0f), .a1 (xffffeeee), .b0 (x33333333), .b1 (xcccccc00));
    nor2b 	m00001110 (.y(x00001110), .an (xfff0fff0), .b  (xffffeeee));
    o22ai 	m00001175 (.y(x00001175), .a0 (x0f0f0f0f), .a1 (xffffffcc), .b0 (xcc00cc00), .b1 (xffffaaaa));
    o22ai 	m00001355 (.y(x00001355), .a0 (x00ff00ff), .a1 (xfffffcfc), .b0 (xcc00cc00), .b1 (xffffaaaa));
    and3 	m00008000 (.y(x00008000), .a  (xf0f0f000), .b  (x88008800), .c  (x0000ffff));
    and3 	m00008880 (.y(x00008880), .a  (x88888888), .b  (xccc0ccc0), .c  (x0000ffff));
    nor2b 	m0000a000 (.y(x0000a000), .an (xa000a000), .b  (xfcfc0000));
    nor2 	m00010005 (.y(x00010005), .a  (xfcfc0000), .b  (xfffafffa));
    o22ai 	m00010031 (.y(x00010031), .a0 (x0f0f0f0f), .a1 (xffffffcc), .b0 (xfcfc0000), .b1 (xffeeffee));
    o22ai 	m00050011 (.y(x00050011), .a0 (x0000ffff), .a1 (xfffafffa), .b0 (xfcfc0000), .b1 (xffeeffee));
    o22ai 	m00050022 (.y(x00050022), .a0 (x0000ffff), .a1 (xfffafffa), .b0 (x55555555), .b1 (xffffffcc));
    o22ai 	m00050300 (.y(x00050300), .a0 (x0000ffff), .a1 (xfffafffa), .b0 (x00ff00ff), .b1 (xfffffcfc));
    o22ai 	m00060006 (.y(x00060006), .a0 (x33333333), .a1 (xfffafffa), .b0 (x55555555), .b1 (xfffcfffc));
    o22ai 	m00070013 (.y(x00070013), .a0 (x0000ffff), .a1 (xfffafffa), .b0 (xf0f0a0a0), .b1 (xffccffcc));
    a31oi 	m0007173f (.y(x0007173f), .a0 (xfcccfccc), .a1 (xeaeaeaea), .a2 (xfffffff0), .b0 (xfff00000));
    a31oi 	m000a022a (.y(x000a022a), .a0 (xfffffcfc), .a1 (xaaa0aaa0), .a2 (xffffffcc), .b0 (x55555555));
    nor2b 	m000a0808 (.y(x000a0808), .an (xaaaa8888), .b  (xfff0f0f0));
    o22ai 	m000aaaab (.y(x000aaaab), .a0 (x55555555), .a1 (xfff00000), .b0 (xfcfccccc), .b1 (xfffffff0));
    nor2 	m000c0e5e (.y(x000c0e5e), .a  (xfff30000), .b  (xf1a1f1a1));
    nor2b 	m000ccc00 (.y(x000ccc00), .an (xcccccc00), .b  (xfff00000));
    o22ai 	m000f023f (.y(x000f023f), .a0 (x55555555), .a1 (xfffffcfc), .b0 (xf0f0c0c0), .b1 (xff00ff00));
    o22ai 	m00113035 (.y(x00113035), .a0 (x0f0f0f0f), .a1 (xf0f0c0c0), .b0 (xccccc0c0), .b1 (xffaaffaa));
    o22ai 	m00130f0f (.y(x00130f0f), .a0 (x0000ffff), .a1 (xffeeffee), .b0 (xfcfc0000), .b1 (xfff0f0f0));
    o22ai 	m00330404 (.y(x00330404), .a0 (x0000ffff), .a1 (xffcc0000), .b0 (x33333333), .b1 (xfffffafa));
    nor4 	m004000c0 (.y(x004000c0), .a  (x88880000), .b  (xf000f000), .c  (x0f0f0f0f), .d  (x33333333));
    o21ai 	m005dccdd (.y(x005dccdd), .a0 (xfff00000), .a1 (x33333333), .b0 (xffaaffaa));
    o22ai 	m007fabff (.y(x007fabff), .a0 (x55555555), .a1 (xfff00000), .b0 (xcc88cc88), .b1 (xff00f000));
    o22ai 	m0100011f (.y(x0100011f), .a0 (x00ff00ff), .a1 (xfefefefe), .b0 (xe0e0e0e0), .b1 (xffffff00));
    o22ai 	m01010003 (.y(x01010003), .a0 (x0000ffff), .a1 (xfefefefe), .b0 (xffaa0000), .b1 (xfffcfffc));
    o22ai 	m01011010 (.y(x01011010), .a0 (x0000ffff), .a1 (xfefefefe), .b0 (x0f0f0f0f), .b1 (xffffeeee));
    o22ai 	m01155fff (.y(x01155fff), .a0 (xeeee0000), .a1 (xf000f000), .b0 (xfafa0000), .b1 (xff00aa00));
    o22ai 	m0133273f (.y(x0133273f), .a0 (x55555555), .a1 (xaaaa8888), .b0 (xccccc0c0), .b1 (xfa00fa00));
    a31oi 	m0137133f (.y(x0137133f), .a0 (xfffff0f0), .a1 (xfafaaaaa), .a2 (xffccffcc), .b0 (xccc0ccc0));
    o22ai 	m01f731f7 (.y(x01f731f7), .a0 (x0f0f0f0f), .a1 (xff00cc00), .b0 (xcc88cc88), .b1 (xfa00fa00));
    nor2b 	m03fc03fc (.y(x03fc03fc), .an (xfffcfffc), .b  (xfc00fc00));
    o22ai 	m04044447 (.y(x04044447), .a0 (x33333333), .a1 (xfafaaaaa), .b0 (xcc88cc88), .b1 (xfffffff0));
    nor4 	m040c0000 (.y(x040c0000), .a  (xc0c00000), .b  (xaa000000), .c  (x33333333), .d  (x0000ffff));
    nor2b 	m05500000 (.y(x05500000), .an (xfff00000), .b  (xfaaafaaa));
    o22ai 	m055f0557 (.y(x055f0557), .a0 (x0000ffff), .a1 (xfff00000), .b0 (xa8a8a8a8), .b1 (xfa00fa00));
    and3 	m08000000 (.y(x08000000), .a  (xfcfc0000), .b  (xaa000000), .c  (x0f0f0f0f));
    nor2b 	m0a000000 (.y(x0a000000), .an (xaa000000), .b  (xf0f00000));
    and3 	m0a080000 (.y(x0a080000), .a  (xaaaa0000), .b  (xffcc0000), .c  (x0f0f0f0f));
    a31oi 	m0abf1bbf (.y(x0abf1bbf), .a0 (xffcccccc), .a1 (x55555555), .a2 (xfff0fff0), .b0 (xa000a000));
    a31oi 	m0b1fafbf (.y(x0b1fafbf), .a0 (xfcccfccc), .a1 (xfff0f0f0), .a2 (x55555555), .b0 (xa0a00000));
    a21oi 	m0cd37660 (.y(x0cd37660), .a0 (xffec8888), .a1 (xf33fffff), .b0 (x00000117));
    and3 	m0e0a0000 (.y(x0e0a0000), .a  (xffaa0000), .b  (xeeee0000), .c  (x0f0f0f0f));
    nor3b 	m0eb6ef2f (.y(x0eb6ef2f), .an (x0ff7ffff), .b  (x01011010), .c  (x004000c0));
    a31oi 	m0f5f0a5f (.y(x0f5f0a5f), .a0 (x55555555), .a1 (xff00ff00), .a2 (x0000ffff), .b0 (xf0a0f0a0));
    a31oi 	m0ff7ffff (.y(x0ff7ffff), .a0 (x88880000), .a1 (x00ff00ff), .a2 (x0f0f0f0f), .b0 (xf0000000));
    nor2b 	m10104040 (.y(x10104040), .an (xf0f0c0c0), .b  (xeeeeaaaa));
    nor2b 	m11004400 (.y(x11004400), .an (xff00cc00), .b  (xeeeeaaaa));
    a21oi 	m11131313 (.y(x11131313), .a0 (xfcfcfcfc), .a1 (xeeeeeeee), .b0 (xaa000000));
    o22ai 	m11771333 (.y(x11771333), .a0 (x0000ffff), .a1 (xeeaaeeaa), .b0 (xa000a000), .b1 (xffcccccc));
    nor2b 	m11aa0000 (.y(x11aa0000), .an (xffaa0000), .b  (xee00ee00));
    a21o 	m12bf5b4f (.y(x12bf5b4f), .a0 (x33ffff0f), .a1 (x0abf1bbf), .b0 (x10104040));
    o22ai 	m131317df (.y(x131317df), .a0 (x33333333), .a1 (xcccccc00), .b0 (xcccc8888), .b1 (xe0e0e0e0));
    o22ai 	m1333131f (.y(x1333131f), .a0 (x0000ffff), .a1 (xffcc0000), .b0 (xcccccc00), .b1 (xe0e0e0e0));
    o22ai 	m135f5fdf (.y(x135f5fdf), .a0 (x33333333), .a1 (xcccccc00), .b0 (xa0a0a0a0), .b1 (xcc000000));
    o22ai 	m13bfbfbf (.y(x13bfbfbf), .a0 (x55555555), .a1 (xff000000), .b0 (xcc000000), .b1 (xe0e0e0e0));
    nor2b 	m15000400 (.y(x15000400), .an (xff00cc00), .b  (xeaeaeaea));
    o22ai 	m151d777f (.y(x151d777f), .a0 (x33333333), .a1 (xccc0ccc0), .b0 (xaaaa8888), .b1 (xc0c00000));
    o22ai 	m15555050 (.y(x15555050), .a0 (x0000ffff), .a1 (xfaaafaaa), .b0 (x0f0f0f0f), .b1 (xeeeeaaaa));
    a31oi 	m169287dc (.y(x169287dc), .a0 (xfcfcf8a0), .a1 (xff7f7f7f), .a2 (xeaefffff), .b0 (x01010003));
    o22ai 	m175f333f (.y(x175f333f), .a0 (x0000ffff), .a1 (xfaaafaaa), .b0 (xa0a00000), .b1 (xccc0ccc0));
    o22ai 	m17ff555f (.y(x17ff555f), .a0 (x0000ffff), .a1 (xfc00fc00), .b0 (xaaa0aaa0), .b1 (xc0c00000));
    a31oi 	m1a10b72b (.y(x1a10b72b), .a0 (xfffff8a0), .a1 (xefefcf8f), .a2 (xf5ff5fff), .b0 (x00000054));
    o22ai 	m1d7f5dff (.y(x1d7f5dff), .a0 (x33333333), .a1 (xf0f0a0a0), .b0 (x88880000), .b1 (xee00ee00));
    a21oi 	m1f7b28d7 (.y(x1f7b28d7), .a0 (x0007173f), .a1 (xffecffa8), .b0 (xe080c000));
    o22ai 	m1f7f55ff (.y(x1f7f55ff), .a0 (x0000ffff), .a1 (xe0e0e0e0), .b0 (x88880000), .b1 (xff00aa00));
    o211ai 	m229616fd (.y(x229616fd), .a0 (xe8e8e800), .a1 (xff010103), .b0 (xdd7fff7f), .c0 (xffffffaa));
    a221oi 	m23369e29 (.y(x23369e29), .a0 (xf003f003), .a1 (x55556666), .b0 (xf0c0f5d5), .b1 (x03fc03fc), .c0 (xcc880000));
    a21oi 	m23853f57 (.y(x23853f57), .a0 (xfefaeca8), .a1 (x557f00ff), .b0 (xc800c000));
    a21boi 	m24cc4461 (.y(x24cc4461), .a0 (x1333131f), .a1 (xfffffffe), .b0n(x37ff5577));
    nor2b 	m2a000000 (.y(x2a000000), .an (xaa000000), .b  (xc0c00000));
    o22ai 	m2aeeaaee (.y(x2aeeaaee), .a0 (x33333333), .a1 (xcc00cc00), .b0 (x55555555), .b1 (xc0c00000));
    o22ai 	m2bffafff (.y(x2bffafff), .a0 (x55555555), .a1 (xc0c00000), .b0 (xcc000000), .b1 (xf000f000));
    o21ai 	m2c6cdf10 (.y(x2c6cdf10), .a0 (xf0a0a0a0), .a1 (x333300cf), .b0 (xdfdf77ff));
    a21oi 	m2ca62526 (.y(x2ca62526), .a0 (xfff8fac8), .a1 (x135f5fdf), .b0 (xc011c011));
    o211ai 	m2d9fb2de (.y(x2d9fb2de), .a0 (xfecccc00), .a1 (xa0a0a1a1), .b0 (xdf77df77), .c0 (xf3f37f7f));
    nor3b 	m2fa5e682 (.y(x2fa5e682), .an (x2fafffff), .b  (x000a0808), .c  (x00001175));
    o21ai 	m2fafffff (.y(x2fafffff), .a0 (xcc000000), .a1 (x55555555), .b0 (xf0f00000));
    nor2b 	m30307000 (.y(x30307000), .an (xf0f0f000), .b  (xcccc8888));
    o22ai 	m3030f1f0 (.y(x3030f1f0), .a0 (x00ff00ff), .a1 (xffffeeee), .b0 (x0f0f0f0f), .b1 (xc0c00000));
    nor2b 	m30c030c0 (.y(x30c030c0), .an (xf0c0f0c0), .b  (xcc00cc00));
    o31a 	m318ab4e1 (.y(x318ab4e1), .a0 (x15000400), .a1 (x30c030c0), .a2 (x000aaaab), .b0 (xbbbbf5f5));
    and3 	m32220000 (.y(x32220000), .a  (xffaa0000), .b  (xfafa0000), .c  (x33333333));
    and3 	m32302020 (.y(x32302020), .a  (xfff0f0f0), .b  (xfafaaaaa), .c  (x33333333));
    a31oi 	m323233fb (.y(x323233fb), .a0 (xffffcccc), .a1 (x55555555), .a2 (x0f0f0f0f), .b0 (xcccccc00));
    a21o 	m326fc4dd (.y(x326fc4dd), .a0 (x005dccdd), .a1 (xc5cfc5df), .b0 (x32220000));
    a31oi 	m333300cf (.y(x333300cf), .a0 (x33333333), .a1 (xfff0fff0), .a2 (x0000ffff), .b0 (xcccccc00));
    a31oi 	m33cfffff (.y(x33cfffff), .a0 (xfcfc0000), .a1 (x00ff00ff), .a2 (x33333333), .b0 (xcc000000));
    a31oi 	m33ffff0f (.y(x33ffff0f), .a0 (xfffff0f0), .a1 (x00ff00ff), .a2 (x0000ffff), .b0 (xcc000000));
    a31oi 	m37303733 (.y(x37303733), .a0 (xffffcccc), .a1 (x00ff00ff), .a2 (x0f0f0f0f), .b0 (xc8c8c8c8));
    o22ai 	m3777053f (.y(x3777053f), .a0 (x0000ffff), .a1 (xcc88cc88), .b0 (xaaaaaa00), .b1 (xf0c0f0c0));
    o22ai 	m37ff5577 (.y(x37ff5577), .a0 (x0000ffff), .a1 (xcc000000), .b0 (xaa88aa88), .b1 (xc0c00000));
    a21o 	m39fe8cff (.y(x39fe8cff), .a0 (xfcfcccff), .a1 (x2bffafff), .b0 (x11aa0000));
    a31oi 	m3c3ffdff (.y(x3c3ffdff), .a0 (xff00aa00), .a1 (x0f0f0f0f), .a2 (x33333333), .b0 (xc0c00000));
    a31oi 	m3cf25843 (.y(x3cf25843), .a0 (x0b1fafbf), .a1 (xfffffffc), .a2 (x77cd77ff), .b0 (xc0008000));
    a21oi 	m3f00ff05 (.y(x3f00ff05), .a0 (x00ff00ff), .a1 (xfffffafa), .b0 (xc0c00000));
    a31oi 	m3f0fffcf (.y(x3f0fffcf), .a0 (xf0f0f0f0), .a1 (x00ff00ff), .a2 (x33333333), .b0 (xc0c00000));
    o22ai 	m3f557fff (.y(x3f557fff), .a0 (x00ff00ff), .a1 (xc000c000), .b0 (xa000a000), .b1 (xffaa0000));
    a31oi 	m3fff2faf (.y(x3fff2faf), .a0 (xfffff0f0), .a1 (x55555555), .a2 (x0000ffff), .b0 (xc000c000));
    nand2 	m3fffffff (.y(x3fffffff), .a  (xc0c00000), .b  (xcc000000));
    nor2b 	m40484048 (.y(x40484048), .an (xc8c8c8c8), .b  (xaaa0aaa0));
    nor2b 	m40c00000 (.y(x40c00000), .an (xc0c00000), .b  (xa000a000));
    a21oi 	m41d5cc5c (.y(x41d5cc5c), .a0 (xf0a0f3a3), .a1 (xbb3333ff), .b0 (x0e0a0000));
    and3b 	m4213e265 (.y(x4213e265), .an (x0000101a), .b  (x4e5feeff), .c  (xf333f377));
    a21oi 	m42e28881 (.y(x42e28881), .a0 (x151d777f), .a1 (xfffffffe), .b0 (xa8000000));
    a31oi 	m4332245f (.y(x4332245f), .a0 (xfcecf8a0), .a1 (xffddddff), .a2 (xbfffffff), .b0 (x00050300));
    a31oi 	m434a8cf5 (.y(x434a8cf5), .a0 (xcccf030f), .a1 (xffffffaa), .a2 (xafa5ffff), .b0 (x30307000));
    a31oi 	m43fecdd2 (.y(x43fecdd2), .a0 (xfeecfaa8), .a1 (xbfbf373f), .a2 (xfd11ffff), .b0 (x00010005));
    a211oi 	m4638af86 (.y(x4638af86), .a0 (x55775071), .a1 (x33cfffff), .b0 (xa8800000), .c0 (x00000008));
    a31oi 	m4e5feeff (.y(x4e5feeff), .a0 (x55555555), .a1 (xff00ff00), .a2 (x33333333), .b0 (xa0a00000));
    and3 	m50004000 (.y(x50004000), .a  (xf0f0f000), .b  (xff00cc00), .c  (x55555555));
    nor3 	m52af6f23 (.y(x52af6f23), .a  (xa8008000), .b  (x05500000), .c  (x000010dc));
    a211o 	m52c516d9 (.y(x52c516d9), .a0 (xfeccfec8), .a1 (x131317df), .b0 (x40c00000), .c0 (x00050011));
    a31oi 	m54eaa319 (.y(x54eaa319), .a0 (xddf7ddf7), .a1 (xfffffeee), .a2 (x01155fff), .b0 (xaa000000));
    nor2b 	m55556666 (.y(x55556666), .an (xffffeeee), .b  (xaaaa8888));
    a31oi 	m55775071 (.y(x55775071), .a0 (x0f0f0f0f), .a1 (xffeeffee), .a2 (x0000ffff), .b0 (xaa88aa88));
    o22ai 	m557f00ff (.y(x557f00ff), .a0 (x0000ffff), .a1 (xaaaa0000), .b0 (xc0c00000), .b1 (xff00ff00));
    o22ai 	m571fff3f (.y(x571fff3f), .a0 (x00ff00ff), .a1 (xaaaa0000), .b0 (xa0a00000), .b1 (xccc0ccc0));
    o22ai 	m57ffff00 (.y(x57ffff00), .a0 (x0000ffff), .a1 (xaa000000), .b0 (x00ff00ff), .b1 (xfcfc0000));
    a31oi 	m5a5f5b5f (.y(x5a5f5b5f), .a0 (xff00cc00), .a1 (x55555555), .a2 (x0f0f0f0f), .b0 (xa0a0a0a0));
    nor2b 	m5aaa5aaa (.y(x5aaa5aaa), .an (xfaaafaaa), .b  (xa000a000));
    a211oi 	m5b847ba9 (.y(x5b847ba9), .a0 (x055f0557), .a1 (xfefafefa), .b0 (xa0008000), .c0 (x00330404));
    a31oi 	m5e9f51e4 (.y(x5e9f51e4), .a0 (xffeeee88), .a1 (xaf7faf7f), .a2 (xf1f1ffff), .b0 (x00000013));
    nor2b 	m5f5ffafa (.y(x5f5ffafa), .an (xfffffafa), .b  (xa0a00000));
    a31oi 	m5fff0faf (.y(x5fff0faf), .a0 (xfffff0f0), .a1 (x55555555), .a2 (x0000ffff), .b0 (xa000a000));
    a211oi 	m6191ae47 (.y(x6191ae47), .a0 (xfeeef8a8), .a1 (x1f7f55ff), .b0 (x88000000), .c0 (x00001110));
    a221oi 	m6a86145f (.y(x6a86145f), .a0 (xdd11cc00), .a1 (x15555050), .b0 (xfff8ffa0), .b1 (x007fabff), .c0 (x80000000));
    or3 	m6ad30f0f (.y(x6ad30f0f), .a  (x2a000000), .b  (x40c00000), .c  (x00130f0f));
    a31oi 	m6d287e63 (.y(x6d287e63), .a0 (x3777053f), .a1 (x5a5f5b5f), .a2 (xfffffffc), .b0 (x80808080));
    a31oi 	m7077f7ff (.y(x7077f7ff), .a0 (xff00cc00), .a1 (xff00aa00), .a2 (x0f0f0f0f), .b0 (x88880000));
    a31oi 	m777717ff (.y(x777717ff), .a0 (xfc00fc00), .a1 (xeaeaeaea), .a2 (x0000ffff), .b0 (x88880000));
    a31oi 	m77cd77ff (.y(x77cd77ff), .a0 (xfafa0000), .a1 (x00ff00ff), .a2 (x33333333), .b0 (x88008800));
    nor2b 	m77fc77fc (.y(x77fc77fc), .an (xfffcfffc), .b  (x88008800));
    a31oi 	m77ff3337 (.y(x77ff3337), .a0 (xfcfccccc), .a1 (xfffafffa), .a2 (x0000ffff), .b0 (x88008800));
    a211o 	m7847e6db (.y(x7847e6db), .a0 (xffcceec8), .a1 (x7077f7ff), .b0 (x08000000), .c0 (x00070013));
    a31oi 	m7c7c7c7d (.y(x7c7c7c7d), .a0 (x0f0f0f0f), .a1 (x33333333), .a2 (xffffffaa), .b0 (x80808080));
    a31oi 	m7ca10f66 (.y(x7ca10f66), .a0 (xfffef888), .a1 (x8fdfffff), .a2 (xf35ff3ff), .b0 (x00001011));
    o22ai 	m7f5f3300 (.y(x7f5f3300), .a0 (x0000ffff), .a1 (xa0a00000), .b0 (x00ff00ff), .b1 (xcc00cc00));
    and2 	m80000000 (.y(x80000000), .a  (xc0c00000), .b  (xa000a000));
    nor3 	m80808080 (.y(x80808080), .a  (x55555555), .b  (x0f0f0f0f), .c  (x33333333));
    o211ai 	m854f7ef5 (.y(x854f7ef5), .a0 (x3030f1f0), .a1 (x5aaa5aaa), .b0 (xfff5f5ff), .c0 (xffff8f0f));
    nor2b 	m88000000 (.y(x88000000), .an (x88880000), .b  (x00ff00ff));
    nor3 	m88008800 (.y(x88008800), .a  (x00ff00ff), .b  (x55555555), .c  (x33333333));
    nor3 	m88880000 (.y(x88880000), .a  (x55555555), .b  (x33333333), .c  (x0000ffff));
    nor2 	m88888888 (.y(x88888888), .a  (x55555555), .b  (x33333333));
    a31oi 	m8ad2e815 (.y(x8ad2e815), .a0 (xffffffea), .a1 (xf5a5ffff), .a2 (x777717ff), .b0 (x040c0000));
    a31oi 	m8b30445b (.y(x8b30445b), .a0 (x77ff3337), .a1 (xffffffec), .a2 (xfccfffff), .b0 (x00008880));
    a21oi 	m8df398a3 (.y(x8df398a3), .a0 (xaa0faf5f), .a1 (x77fc77fc), .b0 (x50004000));
    o22ai 	m8fdfffff (.y(x8fdfffff), .a0 (x33333333), .a1 (x55555555), .b0 (xa0a00000), .b1 (xf0000000));
    a211o 	m96492239 (.y(x96492239), .a0 (xfec8eec8), .a1 (x175f333f), .b0 (x80000000), .c0 (x00010031));
    a21oi 	m9d97aa84 (.y(x9d97aa84), .a0 (xaaaf153f), .a1 (x37303733), .b0 (x40484048));
    and2 	ma0008000 (.y(xa0008000), .a  (xff00cc00), .b  (xa000a000));
    nor3 	ma000a000 (.y(xa000a000), .a  (x00ff00ff), .b  (x55555555), .c  (x0f0f0f0f));
    nor3 	ma0a00000 (.y(xa0a00000), .a  (x55555555), .b  (x0f0f0f0f), .c  (x0000ffff));
    nor2 	ma0a0a0a0 (.y(xa0a0a0a0), .a  (x55555555), .b  (x0f0f0f0f));
    o22ai 	ma0a0a1a1 (.y(xa0a0a1a1), .a0 (x0f0f0f0f), .a1 (x55555555), .b0 (xfcfccccc), .b1 (xfffffafa));
    a31oi 	ma0fb7cd2 (.y(xa0fb7cd2), .a0 (xff05333f), .a1 (x5fff0faf), .a2 (xfffcfffd), .b0 (x00008000));
    o22ai 	ma1b3a5bf (.y(xa1b3a5bf), .a0 (x0f0f0f0f), .a1 (x55555555), .b0 (xccccc0c0), .b1 (xfa00fa00));
    o21ai 	ma4b75f65 (.y(xa4b75f65), .a0 (xfac8a080), .a1 (x0100011f), .b0 (x5f5ffafa));
    and2 	ma8000000 (.y(xa8000000), .a  (xfcfc0000), .b  (xaa000000));
    and3 	ma8008000 (.y(xa8008000), .a  (xfc00fc00), .b  (xff00f000), .c  (xaaaa8888));
    and3 	ma8800000 (.y(xa8800000), .a  (xfff00000), .b  (xffcc0000), .c  (xa8a8a8a8));
    a21oi 	ma8a8a8a8 (.y(xa8a8a8a8), .a0 (x0f0f0f0f), .a1 (x33333333), .b0 (x55555555));
    a21oi 	ma90301b8 (.y(xa90301b8), .a0 (xfaf8fa00), .a1 (x57ffff00), .b0 (x04044447));
    a211oi 	ma9e15289 (.y(xa9e15289), .a0 (xfefea8a0), .a1 (x571fff3f), .b0 (x00060006), .c0 (x00000550));
    nor3 	maa000000 (.y(xaa000000), .a  (x00ff00ff), .b  (x55555555), .c  (x0000ffff));
    o22ai 	maa0faf5f (.y(xaa0faf5f), .a0 (x00ff00ff), .a1 (x55555555), .b0 (xf0f0a0a0), .b1 (xff00f000));
    a21oi 	maa88aa88 (.y(xaa88aa88), .a0 (x00ff00ff), .a1 (x33333333), .b0 (x55555555));
    a21oi 	maaa0aaa0 (.y(xaaa0aaa0), .a0 (x00ff00ff), .a1 (x0f0f0f0f), .b0 (x55555555));
    nor2 	maaaa0000 (.y(xaaaa0000), .a  (x55555555), .b  (x0000ffff));
    a21oi 	maaaa8888 (.y(xaaaa8888), .a0 (x33333333), .a1 (x0000ffff), .b0 (x55555555));
    a21oi 	maaaaa0a0 (.y(xaaaaa0a0), .a0 (x0f0f0f0f), .a1 (x0000ffff), .b0 (x55555555));
    a21oi 	maaaaaa00 (.y(xaaaaaa00), .a0 (x00ff00ff), .a1 (x0000ffff), .b0 (x55555555));
    o22ai 	maaaf153f (.y(xaaaf153f), .a0 (x0000ffff), .a1 (x55555555), .b0 (xf0f0c0c0), .b1 (xff00aa00));
    nand2b 	madffadff (.y(xadffadff), .an (xa8a8a8a8), .b  (xfa00fa00));
    o22ai 	maf7faf7f (.y(xaf7faf7f), .a0 (x00ff00ff), .a1 (x55555555), .b0 (x80808080), .b1 (xf000f000));
    nand2b 	mafa5ffff (.y(xafa5ffff), .an (xaaa0aaa0), .b  (xfafa0000));
    o21a 	mb047c23f (.y(xb047c23f), .a0 (xf0c0c000), .a1 (x000f023f), .b0 (xbb77ffff));
    o22ai 	mb1b1f5f7 (.y(xb1b1f5f7), .a0 (x0f0f0f0f), .a1 (x55555555), .b0 (xaaaaaa00), .b1 (xcccc8888));
    nand2b 	mbb3333ff (.y(xbb3333ff), .an (xaa000000), .b  (xcccccc00));
    o22ai 	mbb77ffff (.y(xbb77ffff), .a0 (x00ff00ff), .a1 (x55555555), .b0 (x88880000), .b1 (xcc000000));
    nand2b 	mbbbbf5f5 (.y(xbbbbf5f5), .an (xaaaaa0a0), .b  (xeeeeaaaa));
    o22ai 	mbfbf373f (.y(xbfbf373f), .a0 (x0000ffff), .a1 (x55555555), .b0 (x88008800), .b1 (xc0c0c0c0));
    nand3 	mbfffffff (.y(xbfffffff), .a  (xc0c00000), .b  (xcc000000), .c  (x55555555));
    and2 	mc0008000 (.y(xc0008000), .a  (xf000f000), .b  (xcccc8888));
    nor3 	mc000c000 (.y(xc000c000), .a  (x00ff00ff), .b  (x0f0f0f0f), .c  (x33333333));
    nand2b 	mc011c011 (.y(xc011c011), .an (xc000c000), .b  (xffeeffee));
    nor3 	mc0c00000 (.y(xc0c00000), .a  (x0f0f0f0f), .b  (x33333333), .c  (x0000ffff));
    nor2 	mc0c0c0c0 (.y(xc0c0c0c0), .a  (x0f0f0f0f), .b  (x33333333));
    o22ai 	mc3c3c3cf (.y(xc3c3c3cf), .a0 (x0f0f0f0f), .a1 (x33333333), .b0 (xcccccc00), .b1 (xf0f0f0f0));
    a21oi 	mc4cf14da (.y(xc4cf14da), .a0 (x3f00ff05), .a1 (xcbffcbff), .b0 (x32302020));
    o22ai 	mc5cfc5df (.y(xc5cfc5df), .a0 (x0f0f0f0f), .a1 (x33333333), .b0 (xf0f0a0a0), .b1 (xfa00fa00));
    o211ai 	mc60b25d3 (.y(xc60b25d3), .a0 (xf8f0c800), .a1 (x0137133f), .b0 (xfffcfeec), .c0 (x3fffffff));
    a21oi 	mc6aca424 (.y(xc6aca424), .a0 (xf8f8c8c8), .a1 (x3f557fff), .b0 (x11131313));
    and2 	mc800c000 (.y(xc800c000), .a  (xff00f000), .b  (xc8c8c8c8));
    a21oi 	mc8c8c8c8 (.y(xc8c8c8c8), .a0 (x55555555), .a1 (x0f0f0f0f), .b0 (x33333333));
    nand2 	mcbea0a80 (.y(xcbea0a80), .a  (xf555f57f), .b  (x3c3ffdff));
    nand2b 	mcbffcbff (.y(xcbffcbff), .an (xc8c8c8c8), .b  (xfc00fc00));
    nor3 	mcc000000 (.y(xcc000000), .a  (x00ff00ff), .b  (x33333333), .c  (x0000ffff));
    nor2 	mcc00cc00 (.y(xcc00cc00), .a  (x00ff00ff), .b  (x33333333));
    nor2b 	mcc880000 (.y(xcc880000), .an (xffaa0000), .b  (x33333333));
    a21oi 	mcc88cc88 (.y(xcc88cc88), .a0 (x00ff00ff), .a1 (x55555555), .b0 (x33333333));
    a21oi 	mccc0ccc0 (.y(xccc0ccc0), .a0 (x00ff00ff), .a1 (x0f0f0f0f), .b0 (x33333333));
    nor2 	mcccc0000 (.y(xcccc0000), .a  (x33333333), .b  (x0000ffff));
    a21oi 	mcccc8888 (.y(xcccc8888), .a0 (x55555555), .a1 (x0000ffff), .b0 (x33333333));
    a21oi 	mccccc0c0 (.y(xccccc0c0), .a0 (x0f0f0f0f), .a1 (x0000ffff), .b0 (x33333333));
    a21oi 	mcccccc00 (.y(xcccccc00), .a0 (x00ff00ff), .a1 (x0000ffff), .b0 (x33333333));
    o22ai 	mcccf030f (.y(xcccf030f), .a0 (x0000ffff), .a1 (x33333333), .b0 (xcc00cc00), .b1 (xfff0f0f0));
    o21ai 	md1f16c3a (.y(xd1f16c3a), .a0 (xeeee8080), .a1 (x00001355), .b0 (x3f0fffcf));
    a21oi 	md2a0de7f (.y(xd2a0de7f), .a0 (xadffadff), .a1 (x7f5f3300), .b0 (x00000080));
    o21ai 	md7997ddd (.y(xd7997ddd), .a0 (xf8008000), .a1 (x11771333), .b0 (x2aeeaaee));
    o22ai 	mdd11cc00 (.y(xdd11cc00), .a0 (x0000ffff), .a1 (xeeee0000), .b0 (x00ff00ff), .b1 (x33333333));
    nand2b 	mdd5555ff (.y(xdd5555ff), .an (xcc000000), .b  (xaaaaaa00));
    o22ai 	mdd7fff7f (.y(xdd7fff7f), .a0 (x00ff00ff), .a1 (x33333333), .b0 (x80808080), .b1 (xaa000000));
    nand2b 	mddf7ddf7 (.y(xddf7ddf7), .an (xccc0ccc0), .b  (xaa88aa88));
    o22ai 	mdf77df77 (.y(xdf77df77), .a0 (x00ff00ff), .a1 (x33333333), .b0 (xa000a000), .b1 (xcc88cc88));
    a21oi 	mdfc11244 (.y(xdfc11244), .a0 (xa1b3a5bf), .a1 (x323233fb), .b0 (x000ccc00));
    o22ai 	mdfdf77ff (.y(xdfdf77ff), .a0 (x0000ffff), .a1 (x33333333), .b0 (x88008800), .b1 (xa0a00000));
    and3 	me080c000 (.y(xe080c000), .a  (xf0f0f000), .b  (xffcccccc), .c  (xeeaaeeaa));
    a21oi 	me0e0e0e0 (.y(xe0e0e0e0), .a0 (x55555555), .a1 (x33333333), .b0 (x0f0f0f0f));
    nand3b 	me2cda26e (.y(xe2cda26e), .an (x00050022), .b  (x1d7f5dff), .c  (xffb3ffb3));
    a31oi 	me3ab5bd2 (.y(xe3ab5bd2), .a0 (x7c7c7c7d), .a1 (xdd5555ff), .a2 (x3fff2faf), .b0 (x0000a000));
    a21oi 	me8133bb7 (.y(xe8133bb7), .a0 (xffecece8), .a1 (x17ff555f), .b0 (x00008000));
    and3 	me8e8e800 (.y(xe8e8e800), .a  (xfcfcfcfc), .b  (xeaeaeaea), .c  (xffffff00));
    o21ai 	meaeaeaea (.y(xeaeaeaea), .a0 (x0f0f0f0f), .a1 (x33333333), .b0 (x55555555));
    nand2b 	meaefffff (.y(xeaefffff), .an (xeaeaeaea), .b  (xfff00000));
    a21oi 	mee00ee00 (.y(xee00ee00), .a0 (x55555555), .a1 (x33333333), .b0 (x00ff00ff));
    o21ai 	meeaaeeaa (.y(xeeaaeeaa), .a0 (x00ff00ff), .a1 (x33333333), .b0 (x55555555));
    a21oi 	meecc98e2 (.y(xeecc98e2), .a0 (x0133273f), .a1 (xffffffdd), .b0 (x11004400));
    a21oi 	meeee0000 (.y(xeeee0000), .a0 (x55555555), .a1 (x33333333), .b0 (x0000ffff));
    or2 	meeee8080 (.y(xeeee8080), .a  (xeeee0000), .b  (x80808080));
    o21ai 	meeeeaaaa (.y(xeeeeaaaa), .a0 (x33333333), .a1 (x0000ffff), .b0 (x55555555));
    nand2 	meeeeeeee (.y(xeeeeeeee), .a  (x55555555), .b  (x33333333));
    a21oi 	mef715dd5 (.y(xef715dd5), .a0 (xfccca000), .a1 (x13bfbfbf), .b0 (x000a022a));
    or3 	mefefcf8f (.y(xefefcf8f), .a  (xeeee0000), .b  (xcc88cc88), .c  (x0f0f0f0f));
    nor3 	mf0000000 (.y(xf0000000), .a  (x00ff00ff), .b  (x0f0f0f0f), .c  (x0000ffff));
    nor2 	mf000f000 (.y(xf000f000), .a  (x00ff00ff), .b  (x0f0f0f0f));
    nand2b 	mf003f003 (.y(xf003f003), .an (xf000f000), .b  (xfffcfffc));
    nor2b 	mf0a0a0a0 (.y(xf0a0a0a0), .an (xffaaaaaa), .b  (x0f0f0f0f));
    a21oi 	mf0a0f0a0 (.y(xf0a0f0a0), .a0 (x00ff00ff), .a1 (x55555555), .b0 (x0f0f0f0f));
    nand2b 	mf0a0f3a3 (.y(xf0a0f3a3), .an (xf0a0f0a0), .b  (xfffffcfc));
    and2 	mf0c0c000 (.y(xf0c0c000), .a  (xf0f0f000), .b  (xffcccccc));
    a21oi 	mf0c0f0c0 (.y(xf0c0f0c0), .a0 (x00ff00ff), .a1 (x33333333), .b0 (x0f0f0f0f));
    nand2b 	mf0c0f5d5 (.y(xf0c0f5d5), .an (xf0c0f0c0), .b  (xffffaaaa));
    nor2 	mf0f00000 (.y(xf0f00000), .a  (x0f0f0f0f), .b  (x0000ffff));
    a21oi 	mf0f0a0a0 (.y(xf0f0a0a0), .a0 (x55555555), .a1 (x0000ffff), .b0 (x0f0f0f0f));
    a21oi 	mf0f0c0c0 (.y(xf0f0c0c0), .a0 (x33333333), .a1 (x0000ffff), .b0 (x0f0f0f0f));
    a21oi 	mf0f0f000 (.y(xf0f0f000), .a0 (x00ff00ff), .a1 (x0000ffff), .b0 (x0f0f0f0f));
    inv 	mf0f0f0f0 (.y(xf0f0f0f0), .a  (x0f0f0f0f));
    and3b 	mf12405c2 (.y(xf12405c2), .an (x00113035), .b  (xf1f5f5f7), .c  (xff3f05ff));
    nand2b 	mf1a1f1a1 (.y(xf1a1f1a1), .an (xf0a0f0a0), .b  (xfefefefe));
    nand2 	mf1f1ffff (.y(xf1f1ffff), .a  (xeeee0000), .b  (x0f0f0f0f));
    nand4 	mf1f5f5f7 (.y(xf1f5f5f7), .a  (xeeeeaaaa), .b  (xffaaaaaa), .c  (x0f0f0f0f), .d  (xffffffcc));
    o22ai 	mf333f377 (.y(xf333f377), .a0 (x00ff00ff), .a1 (x0f0f0f0f), .b0 (xcc00cc00), .b1 (xcccc8888));
    o22ai 	mf33fffff (.y(xf33fffff), .a0 (x00ff00ff), .a1 (x0f0f0f0f), .b0 (xc0c00000), .b1 (xcc000000));
    o22ai 	mf35ff3ff (.y(xf35ff3ff), .a0 (x00ff00ff), .a1 (x0f0f0f0f), .b0 (xa0a00000), .b1 (xcc00cc00));
    o22ai 	mf3f37f7f (.y(xf3f37f7f), .a0 (x0000ffff), .a1 (x0f0f0f0f), .b0 (x80808080), .b1 (xfcfc0000));
    a21oi 	mf446ce08 (.y(xf446ce08), .a0 (x01f731f7), .a1 (xb1b1f5f7), .b0 (x0a080000));
    a21oi 	mf4bcfdb0 (.y(xf4bcfdb0), .a0 (x0f5f0a5f), .a1 (xc3c3c3cf), .b0 (x0a000000));
    o22ai 	mf555f57f (.y(xf555f57f), .a0 (x00ff00ff), .a1 (x0f0f0f0f), .b0 (x80808080), .b1 (xaaaaaa00));
    nand2b 	mf5a5ffff (.y(xf5a5ffff), .an (xf0a0f0a0), .b  (xfafa0000));
    o22ai 	mf5ff5fff (.y(xf5ff5fff), .a0 (x0000ffff), .a1 (x0f0f0f0f), .b0 (xa000a000), .b1 (xaa000000));
    and3 	mf8008000 (.y(xf8008000), .a  (xff00f000), .b  (xfcfccccc), .c  (xfafaaaaa));
    or3 	mf8f0c800 (.y(xf8f0c800), .a  (xf0f00000), .b  (x88008800), .c  (xc000c000));
    and2 	mf8f8c8c8 (.y(xf8f8c8c8), .a  (xfcfccccc), .b  (xfafafafa));
    a21oi 	mfa00fa00 (.y(xfa00fa00), .a0 (x55555555), .a1 (x0f0f0f0f), .b0 (x00ff00ff));
    o21ai 	mfaaafaaa (.y(xfaaafaaa), .a0 (x00ff00ff), .a1 (x0f0f0f0f), .b0 (x55555555));
    and3 	mfac8a080 (.y(xfac8a080), .a  (xfffff0f0), .b  (xfafaaaaa), .c  (xffccffcc));
    and3 	mfaf8fa00 (.y(xfaf8fa00), .a  (xfafafafa), .b  (xffffff00), .c  (xfffcfffc));
    a21oi 	mfafa0000 (.y(xfafa0000), .a0 (x55555555), .a1 (x0f0f0f0f), .b0 (x0000ffff));
    o21ai 	mfafaaaaa (.y(xfafaaaaa), .a0 (x0f0f0f0f), .a1 (x0000ffff), .b0 (x55555555));
    nand2 	mfafafafa (.y(xfafafafa), .a  (x55555555), .b  (x0f0f0f0f));
    a21oi 	mfc00fc00 (.y(xfc00fc00), .a0 (x0f0f0f0f), .a1 (x33333333), .b0 (x00ff00ff));
    or3 	mfccca000 (.y(xfccca000), .a  (xcccc0000), .b  (xa000a000), .c  (xf0000000));
    o21ai 	mfcccfccc (.y(xfcccfccc), .a0 (x00ff00ff), .a1 (x0f0f0f0f), .b0 (x33333333));
    nand2b 	mfccfffff (.y(xfccfffff), .an (xfcccfccc), .b  (xfff00000));
    or3 	mfcecf8a0 (.y(xfcecf8a0), .a  (xcccc0000), .b  (x88008800), .c  (xf0a0f0a0));
    a21oi 	mfcfc0000 (.y(xfcfc0000), .a0 (x0f0f0f0f), .a1 (x33333333), .b0 (x0000ffff));
    o21ai 	mfcfccccc (.y(xfcfccccc), .a0 (x0f0f0f0f), .a1 (x0000ffff), .b0 (x33333333));
    nand2b 	mfcfcccff (.y(xfcfcccff), .an (xfcfccccc), .b  (xffffff00));
    or3 	mfcfcf8a0 (.y(xfcfcf8a0), .a  (xfcfc0000), .b  (x88008800), .c  (xf0a0f0a0));
    nand2 	mfcfcfcfc (.y(xfcfcfcfc), .a  (x0f0f0f0f), .b  (x33333333));
    nand2b 	mfd11ffff (.y(xfd11ffff), .an (xfc00fc00), .b  (xeeee0000));
    or3 	mfec8eec8 (.y(xfec8eec8), .a  (xf0000000), .b  (xccc0ccc0), .c  (xaa88aa88));
    and3 	mfecccc00 (.y(xfecccc00), .a  (xffcccccc), .b  (xfefefefe), .c  (xffffff00));
    or3 	mfeccfec8 (.y(xfeccfec8), .a  (xfc00fc00), .b  (xccccc0c0), .c  (xaa88aa88));
    or3 	mfeecfaa8 (.y(xfeecfaa8), .a  (xf000f000), .b  (xcccc8888), .c  (xaaa0aaa0));
    or3 	mfeeef8a8 (.y(xfeeef8a8), .a  (xf000f000), .b  (xeeee0000), .c  (xa8a8a8a8));
    or3 	mfefaeca8 (.y(xfefaeca8), .a  (xcc00cc00), .b  (xfafa0000), .c  (xa8a8a8a8));
    nand2b 	mfefafefa (.y(xfefafefa), .an (xeeaaeeaa), .b  (x0f0f0f0f));
    or3 	mfefea8a0 (.y(xfefea8a0), .a  (xfcfc0000), .b  (x88008800), .c  (xaaaaa0a0));
    nand3 	mfefefefe (.y(xfefefefe), .a  (x55555555), .b  (x0f0f0f0f), .c  (x33333333));
    nor2 	mff000000 (.y(xff000000), .a  (x00ff00ff), .b  (x0000ffff));
    a21oi 	mff00aa00 (.y(xff00aa00), .a0 (x55555555), .a1 (x0000ffff), .b0 (x00ff00ff));
    a21oi 	mff00cc00 (.y(xff00cc00), .a0 (x33333333), .a1 (x0000ffff), .b0 (x00ff00ff));
    a21oi 	mff00f000 (.y(xff00f000), .a0 (x0f0f0f0f), .a1 (x0000ffff), .b0 (x00ff00ff));
    inv 	mff00ff00 (.y(xff00ff00), .a  (x00ff00ff));
    o22ai 	mff010103 (.y(xff010103), .a0 (x0000ffff), .a1 (x00ff00ff), .b0 (xaaaaaa00), .b1 (xfcfcfcfc));
    o22ai 	mff05333f (.y(xff05333f), .a0 (x0000ffff), .a1 (x00ff00ff), .b0 (xccc0ccc0), .b1 (xfafa0000));
    o22ai 	mff3f05ff (.y(xff3f05ff), .a0 (x0000ffff), .a1 (x00ff00ff), .b0 (xc0c00000), .b1 (xfa00fa00));
    nand2b 	mff7f7f7f (.y(xff7f7f7f), .an (xcc000000), .b  (x80808080));
    a21oi 	mffaa0000 (.y(xffaa0000), .a0 (x00ff00ff), .a1 (x55555555), .b0 (x0000ffff));
    o21ai 	mffaaaaaa (.y(xffaaaaaa), .a0 (x00ff00ff), .a1 (x0000ffff), .b0 (x55555555));
    nand2 	mffaaffaa (.y(xffaaffaa), .a  (x00ff00ff), .b  (x55555555));
    or3 	mffb3ffb3 (.y(xffb3ffb3), .a  (xcc00cc00), .b  (x80808080), .c  (x33333333));
    a21oi 	mffcc0000 (.y(xffcc0000), .a0 (x00ff00ff), .a1 (x33333333), .b0 (x0000ffff));
    o21ai 	mffcccccc (.y(xffcccccc), .a0 (x00ff00ff), .a1 (x0000ffff), .b0 (x33333333));
    or3 	mffcceec8 (.y(xffcceec8), .a  (xff00cc00), .b  (xccccc0c0), .c  (xaa88aa88));
    nand2 	mffccffcc (.y(xffccffcc), .a  (x00ff00ff), .b  (x33333333));
    nand2b 	mffddddff (.y(xffddddff), .an (xffcccccc), .b  (xaaaaaa00));
    or3 	mffec8888 (.y(xffec8888), .a  (xff000000), .b  (xa0a00000), .c  (xcccc8888));
    or3 	mffecece8 (.y(xffecece8), .a  (xff00cc00), .b  (xcccc8888), .c  (xe0e0e0e0));
    and3 	mffecffa8 (.y(xffecffa8), .a  (xffffffaa), .b  (xffeeffee), .c  (xfffcfffc));
    or3 	mffeeee88 (.y(xffeeee88), .a  (xffaa0000), .b  (xcccccc00), .c  (xaa88aa88));
    nand3 	mffeeffee (.y(xffeeffee), .a  (x00ff00ff), .b  (x55555555), .c  (x33333333));
    a21oi 	mfff00000 (.y(xfff00000), .a0 (x00ff00ff), .a1 (x0f0f0f0f), .b0 (x0000ffff));
    o21ai 	mfff0f0f0 (.y(xfff0f0f0), .a0 (x00ff00ff), .a1 (x0000ffff), .b0 (x0f0f0f0f));
    nand2 	mfff0fff0 (.y(xfff0fff0), .a  (x00ff00ff), .b  (x0f0f0f0f));
    a31oi 	mfff30000 (.y(xfff30000), .a0 (xfcfc0000), .a1 (x00ff00ff), .a2 (x0f0f0f0f), .b0 (x0000ffff));
    nand2b 	mfff5f5ff (.y(xfff5f5ff), .an (xfff0f0f0), .b  (xaaaaaa00));
    or3 	mfff8fac8 (.y(xfff8fac8), .a  (xfff00000), .b  (xf0c0f0c0), .c  (xaa88aa88));
    or3 	mfff8ffa0 (.y(xfff8ffa0), .a  (x88880000), .b  (xf0f0a0a0), .c  (xff00ff00));
    nand3 	mfffafffa (.y(xfffafffa), .a  (x00ff00ff), .b  (x55555555), .c  (x0f0f0f0f));
    or3 	mfffcfeec (.y(xfffcfeec), .a  (xf0f0f000), .b  (xffcccccc), .c  (xaaa0aaa0));
    nand3 	mfffcfffc (.y(xfffcfffc), .a  (x00ff00ff), .b  (x0f0f0f0f), .c  (x33333333));
    nand2b 	mfffcfffd (.y(xfffcfffd), .an (xfffcfffc), .b  (xffffaaaa));
    or3 	mfffef888 (.y(xfffef888), .a  (xfcfc0000), .b  (xff00f000), .c  (xaaaa8888));
    inv 	mffff0000 (.y(xffff0000), .a  (x0000ffff));
    or3 	mffff8f0f (.y(xffff8f0f), .a  (xfcfc0000), .b  (x88008800), .c  (x0f0f0f0f));
    nand2 	mffffaaaa (.y(xffffaaaa), .a  (x55555555), .b  (x0000ffff));
    nand2 	mffffcccc (.y(xffffcccc), .a  (x33333333), .b  (x0000ffff));
    nand3 	mffffeeee (.y(xffffeeee), .a  (x55555555), .b  (x33333333), .c  (x0000ffff));
    nand2 	mfffff0f0 (.y(xfffff0f0), .a  (x0f0f0f0f), .b  (x0000ffff));
    or3 	mfffff8a0 (.y(xfffff8a0), .a  (xffff0000), .b  (x88008800), .c  (xf0a0f0a0));
    nand3 	mfffffafa (.y(xfffffafa), .a  (x55555555), .b  (x0f0f0f0f), .c  (x0000ffff));
    nand3 	mfffffcfc (.y(xfffffcfc), .a  (x0f0f0f0f), .b  (x33333333), .c  (x0000ffff));
    or2 	mfffffeee (.y(xfffffeee), .a  (xf0f0f000), .b  (xffffeeee));
    nand2 	mffffff00 (.y(xffffff00), .a  (x00ff00ff), .b  (x0000ffff));
    nand3 	mffffffaa (.y(xffffffaa), .a  (x00ff00ff), .b  (x55555555), .c  (x0000ffff));
    nand3 	mffffffcc (.y(xffffffcc), .a  (x00ff00ff), .b  (x33333333), .c  (x0000ffff));
    nand2b 	mffffffdd (.y(xffffffdd), .an (xffffffcc), .b  (xeeeeaaaa));
    or2 	mffffffea (.y(xffffffea), .a  (xf0f0c0c0), .b  (xffffffaa));
    or2 	mffffffec (.y(xffffffec), .a  (xf0f0a0a0), .b  (xffffffcc));
    nand3 	mfffffff0 (.y(xfffffff0), .a  (x00ff00ff), .b  (x0f0f0f0f), .c  (x0000ffff));
    nand2b 	mfffffffc (.y(xfffffffc), .an (xfffffcfc), .b  (x00ff00ff));
    or2 	mfffffffe (.y(xfffffffe), .a  (xffffcccc), .b  (xfffafffa));

    a22oi   m0a (.y(x0a), .a0(x80), .a1(x52af6f23), .b0(x40), .b1(x4332245f));
    a22oi   m0b (.y(x0b), .a0(x20), .a1(x000c0e5e), .b0(x10), .b1(x229616fd));
    a22oi   m0c (.y(x0c), .a0(x08), .a1(x7ca10f66), .b0(x04), .b1(xdfc11244));
    a22oi   m0d (.y(x0d), .a0(x02), .a1(xd7997ddd), .b0(x01), .b1(x326fc4dd));
    nand4   m0  (.y(x0), .a(x0a), .b(x0b), .c(x0c), .d(x0d));

    a22oi   m1a (.y(x1a), .a0(x80), .a1(xa4b75f65), .b0(x40), .b1(x5e9f51e4));
    a22oi   m1b (.y(x1b), .a0(x20), .a1(xa90301b8), .b0(x10), .b1(x23853f57));
    a22oi   m1c (.y(x1c), .a0(x08), .a1(x8df398a3), .b0(x04), .b1(xa0fb7cd2));
    a22oi   m1d (.y(x1d), .a0(x02), .a1(x96492239), .b0(x01), .b1(x2c6cdf10));
    nand4   m1  (.y(x1), .a(x1a), .b(x1b), .c(x1c), .d(x1d));

    a22oi   m2a (.y(x2a), .a0(x80), .a1(x169287dc), .b0(x40), .b1(xa9e15289));
    a22oi   m2b (.y(x2b), .a0(x20), .a1(x39fe8cff), .b0(x10), .b1(x0cd37660));
    a22oi   m2c (.y(x2c), .a0(x08), .a1(x0eb6ef2f), .b0(x04), .b1(x8ad2e815));
    a22oi   m2d (.y(x2d), .a0(x02), .a1(xc60b25d3), .b0(x01), .b1(x1a10b72b));
    nand4   m2  (.y(x2), .a(x2a), .b(x2b), .c(x2c), .d(x2d));

    a22oi   m3a (.y(x3a), .a0(x80), .a1(x6191ae47), .b0(x40), .b1(x41d5cc5c));
    a22oi   m3b (.y(x3b), .a0(x20), .a1(x4638af86), .b0(x10), .b1(x6d287e63));
    a22oi   m3c (.y(x3c), .a0(x08), .a1(x8b30445b), .b0(x04), .b1(x2d9fb2de));
    a22oi   m3d (.y(x3d), .a0(x02), .a1(xe8133bb7), .b0(x01), .b1(x3cf25843));
    nand4   m3  (.y(x3), .a(x3a), .b(x3b), .c(x3c), .d(x3d));

    a22oi   m4a (.y(x4a), .a0(x80), .a1(x9d97aa84), .b0(x40), .b1(xf12405c2));
    a22oi   m4b (.y(x4b), .a0(x20), .a1(xe3ab5bd2), .b0(x10), .b1(xc6aca424));
    a22oi   m4c (.y(x4c), .a0(x08), .a1(xe2cda26e), .b0(x04), .b1(x7847e6db));
    a22oi   m4d (.y(x4d), .a0(x02), .a1(xd1f16c3a), .b0(x01), .b1(x23369e29));
    nand4   m4  (.y(x4), .a(x4a), .b(x4b), .c(x4c), .d(x4d));

    a22oi   m5a (.y(x5a), .a0(x80), .a1(x2fa5e682), .b0(x40), .b1(x5b847ba9));
    a22oi   m5b (.y(x5b), .a0(x20), .a1(xf446ce08), .b0(x10), .b1(x24cc4461));
    a22oi   m5c (.y(x5c), .a0(x08), .a1(x854f7ef5), .b0(x04), .b1(x54eaa319));
    a22oi   m5d (.y(x5d), .a0(x02), .a1(x318ab4e1), .b0(x01), .b1(xef715dd5));
    nand4   m5  (.y(x5), .a(x5a), .b(x5b), .c(x5c), .d(x5d));

    a22oi   m6a (.y(x6a), .a0(x80), .a1(xb047c23f), .b0(x40), .b1(xc4cf14da));
    a22oi   m6b (.y(x6b), .a0(x20), .a1(xf4bcfdb0), .b0(x10), .b1(x42e28881));
    a22oi   m6c (.y(x6c), .a0(x08), .a1(x1f7b28d7), .b0(x04), .b1(xd2a0de7f));
    a22oi   m6d (.y(x6d), .a0(x02), .a1(x4213e265), .b0(x01), .b1(x52c516d9));
    nand4   m6  (.y(x6), .a(x6a), .b(x6b), .c(x6c), .d(x6d));

    a22oi   m7a (.y(x7a), .a0(x80), .a1(x12bf5b4f), .b0(x40), .b1(x2ca62526));
    a22oi   m7b (.y(x7b), .a0(x20), .a1(x6ad30f0f), .b0(x10), .b1(xeecc98e2));
    a22oi   m7c (.y(x7c), .a0(x08), .a1(x43fecdd2), .b0(x04), .b1(x434a8cf5));
    a22oi   m7d (.y(x7d), .a0(x02), .a1(x6a86145f), .b0(x01), .b1(xcbea0a80));
    nand4   m7  (.y(x7), .a(x7a), .b(x7b), .c(x7c), .d(x7d));

    assign y[7] = x7;
    assign y[6] = x6;
    assign y[5] = x5;
    assign y[4] = x4;
    assign y[3] = x3;
    assign y[2] = x2;
    assign y[1] = x1;
    assign y[0] = x0;

    always @(posedge clk)
    begin
        cy[7] <= x7;
        cy[6] <= x6;
        cy[5] <= x5;
        cy[4] <= x4;
        cy[3] <= x3;
        cy[2] <= x2;
        cy[1] <= x1;
        cy[0] <= x0;
    end

endmodule
