module byte_transmitter_formal ();
endmodule
