module i2c_periph_formal ();

endmodule
