/*
 * Copyright (c) 2024 Your Name
 * SPDX-License-Identifier: Apache-2.0
 */

`default_nettype none

module tt_um_sign_addsub (
    input  wire [7:0] ui_in,    // Dedicated inputs
    output wire [7:0] uo_out,   // Dedicated outputs
    input  wire [7:0] uio_in,   // IOs: Input path
    output wire [7:0] uio_out,  // IOs: Output path
    output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // always 1 when the design is powered, so you can ignore it
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);


 // assign uo_out  = ui_in + uio_in;  // Example: ou_out is the sum of ui_in and uio_in
  signed_addsub_4 A1 (	.a(ui_in[3:0]),
						.b(ui_in[7:4]), 
						.res_signed(uo_out[3:0]),
						.sign(uio_in[1:0]));

   // All output pins must be assigned. If not used, assign to 0.
   assign uo_out[7:4] = 0;
   assign uio_out = 0;

   // List all unused inputs to prevent warnings
  // assign uio_in[7:2] = 0;
  assign uio_oe  = 0;
  wire _unused = &{ena, clk, rst_n, uio_in[7:2], 1'b0};

endmodule

//-----------------------------------------------------------------------------------------------------------------------------------------------------	

