`define SINE_IN_BITS  8
`define SINE_OUT_BITS 8
