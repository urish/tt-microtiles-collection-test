module keccakf1600_statepermutate_tb;
  reg clk;
  reg rstn;
  reg [64*24-1:0] din;
  wire [64*24-1:0] dout;

  keccakf1600_statepermutate uut (
    .clk(clk),
    .rstn(rstn),
    .din(din),
    .dout(dout)
  );

  always #5 clk = ~clk; 

  initial begin
    clk = 0;
    rstn = 0;
    din = {
      64'h0000000000000001,
      64'h0000000000000002,
      64'h0000000000000003,
      64'h0000000000000004,
      64'h0000000000000005,
      64'h0000000000000006,
      64'h0000000000000007,
      64'h0000000000000008,
      64'h0000000000000009,
      64'h000000000000000A,
      64'h000000000000000B,
      64'h000000000000000C,
      64'h000000000000000D,
      64'h000000000000000E,
      64'h000000000000000F,
      64'h0000000000000010,
      64'h0000000000000011,
      64'h0000000000000012,
      64'h0000000000000013,
      64'h0000000000000014,
      64'h0000000000000015,
      64'h0000000000000016,
      64'h0000000000000017,
      64'h0000000000000018,
      64'h0000000000000019
    };


    #10 rstn = 1;  

    #1000; 

    $finish; 
  end

endmodule
