module sky130_fd_sc_hd_dlygate4sd3_1 (
    input A,
    output reg X
);
    sky130_fd_sc_hd__dlygate4sd3_1 i (
        .A(A),
        .X(X)
    );
endmodule
