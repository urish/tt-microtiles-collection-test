//
// SPDX-FileCopyrightText: Copyright 2023 Darryl Miles
// SPDX-License-Identifier: Apache2.0
//

`define UIO_OE_INPUT   1'b0
`define UIO_OE_OUTPUT  1'b1
