/*
 * Copyright (c) 2024 Uri Shaked
 * SPDX-License-Identifier: Apache-2.0
 */

module glyph_2 (
    input wire [5:0] x,
    input wire [5:0] y,
    output wire pixel
);

  reg [7:0] mem[511:0];
  initial begin
    mem[0] = 8'h00;
    mem[1] = 8'h00;
    mem[2] = 8'h00;
    mem[3] = 8'h00;
    mem[4] = 8'h00;
    mem[5] = 8'h00;
    mem[6] = 8'h00;
    mem[7] = 8'h00;
    mem[8] = 8'h00;
    mem[9] = 8'h00;
    mem[10] = 8'h00;
    mem[11] = 8'h00;
    mem[12] = 8'h00;
    mem[13] = 8'h00;
    mem[14] = 8'h00;
    mem[15] = 8'h00;
    mem[16] = 8'h00;
    mem[17] = 8'h00;
    mem[18] = 8'h00;
    mem[19] = 8'h00;
    mem[20] = 8'h00;
    mem[21] = 8'h00;
    mem[22] = 8'h00;
    mem[23] = 8'h00;
    mem[24] = 8'h00;
    mem[25] = 8'h00;
    mem[26] = 8'h00;
    mem[27] = 8'h00;
    mem[28] = 8'h00;
    mem[29] = 8'h00;
    mem[30] = 8'h00;
    mem[31] = 8'h00;
    mem[32] = 8'h00;
    mem[33] = 8'h00;
    mem[34] = 8'h00;
    mem[35] = 8'h00;
    mem[36] = 8'h00;
    mem[37] = 8'h00;
    mem[38] = 8'h00;
    mem[39] = 8'h00;
    mem[40] = 8'h00;
    mem[41] = 8'h00;
    mem[42] = 8'h00;
    mem[43] = 8'h00;
    mem[44] = 8'h00;
    mem[45] = 8'h00;
    mem[46] = 8'h00;
    mem[47] = 8'h00;
    mem[48] = 8'h00;
    mem[49] = 8'h00;
    mem[50] = 8'h00;
    mem[51] = 8'h00;
    mem[52] = 8'h00;
    mem[53] = 8'h00;
    mem[54] = 8'h00;
    mem[55] = 8'h00;
    mem[56] = 8'h00;
    mem[57] = 8'h00;
    mem[58] = 8'h00;
    mem[59] = 8'h00;
    mem[60] = 8'h00;
    mem[61] = 8'h00;
    mem[62] = 8'h00;
    mem[63] = 8'h00;
    mem[64] = 8'h00;
    mem[65] = 8'h00;
    mem[66] = 8'h00;
    mem[67] = 8'h00;
    mem[68] = 8'h00;
    mem[69] = 8'h00;
    mem[70] = 8'h00;
    mem[71] = 8'h00;
    mem[72] = 8'h00;
    mem[73] = 8'h00;
    mem[74] = 8'h00;
    mem[75] = 8'h00;
    mem[76] = 8'h00;
    mem[77] = 8'h00;
    mem[78] = 8'h00;
    mem[79] = 8'h00;
    mem[80] = 8'h00;
    mem[81] = 8'h00;
    mem[82] = 8'h00;
    mem[83] = 8'h00;
    mem[84] = 8'h00;
    mem[85] = 8'h00;
    mem[86] = 8'h00;
    mem[87] = 8'h00;
    mem[88] = 8'h00;
    mem[89] = 8'h00;
    mem[90] = 8'h00;
    mem[91] = 8'h00;
    mem[92] = 8'h00;
    mem[93] = 8'h00;
    mem[94] = 8'h00;
    mem[95] = 8'h00;
    mem[96] = 8'h00;
    mem[97] = 8'h00;
    mem[98] = 8'h00;
    mem[99] = 8'h00;
    mem[100] = 8'h00;
    mem[101] = 8'h00;
    mem[102] = 8'h00;
    mem[103] = 8'h00;
    mem[104] = 8'h00;
    mem[105] = 8'h00;
    mem[106] = 8'h00;
    mem[107] = 8'h00;
    mem[108] = 8'h00;
    mem[109] = 8'h00;
    mem[110] = 8'h00;
    mem[111] = 8'h00;
    mem[112] = 8'h00;
    mem[113] = 8'h00;
    mem[114] = 8'h00;
    mem[115] = 8'h00;
    mem[116] = 8'h00;
    mem[117] = 8'h00;
    mem[118] = 8'h00;
    mem[119] = 8'h00;
    mem[120] = 8'h00;
    mem[121] = 8'h00;
    mem[122] = 8'h00;
    mem[123] = 8'h00;
    mem[124] = 8'h00;
    mem[125] = 8'h00;
    mem[126] = 8'h00;
    mem[127] = 8'h00;
    mem[128] = 8'h00;
    mem[129] = 8'h00;
    mem[130] = 8'h00;
    mem[131] = 8'h00;
    mem[132] = 8'h00;
    mem[133] = 8'h00;
    mem[134] = 8'h00;
    mem[135] = 8'h00;
    mem[136] = 8'h00;
    mem[137] = 8'h00;
    mem[138] = 8'h00;
    mem[139] = 8'hf0;
    mem[140] = 8'h3f;
    mem[141] = 8'h00;
    mem[142] = 8'h00;
    mem[143] = 8'h00;
    mem[144] = 8'h00;
    mem[145] = 8'h00;
    mem[146] = 8'h00;
    mem[147] = 8'hfc;
    mem[148] = 8'hff;
    mem[149] = 8'h00;
    mem[150] = 8'h00;
    mem[151] = 8'h00;
    mem[152] = 8'h00;
    mem[153] = 8'h00;
    mem[154] = 8'h00;
    mem[155] = 8'hfe;
    mem[156] = 8'hff;
    mem[157] = 8'h01;
    mem[158] = 8'h00;
    mem[159] = 8'h00;
    mem[160] = 8'h00;
    mem[161] = 8'h00;
    mem[162] = 8'h00;
    mem[163] = 8'h1f;
    mem[164] = 8'hf0;
    mem[165] = 8'h03;
    mem[166] = 8'h00;
    mem[167] = 8'h00;
    mem[168] = 8'h00;
    mem[169] = 8'h00;
    mem[170] = 8'h00;
    mem[171] = 8'h0f;
    mem[172] = 8'he0;
    mem[173] = 8'h07;
    mem[174] = 8'h00;
    mem[175] = 8'h00;
    mem[176] = 8'h00;
    mem[177] = 8'h00;
    mem[178] = 8'h80;
    mem[179] = 8'h07;
    mem[180] = 8'hc0;
    mem[181] = 8'h07;
    mem[182] = 8'h00;
    mem[183] = 8'h00;
    mem[184] = 8'h00;
    mem[185] = 8'h00;
    mem[186] = 8'h80;
    mem[187] = 8'h07;
    mem[188] = 8'h80;
    mem[189] = 8'h07;
    mem[190] = 8'h00;
    mem[191] = 8'h00;
    mem[192] = 8'h00;
    mem[193] = 8'h00;
    mem[194] = 8'hc0;
    mem[195] = 8'h07;
    mem[196] = 8'h80;
    mem[197] = 8'h07;
    mem[198] = 8'h00;
    mem[199] = 8'h00;
    mem[200] = 8'h00;
    mem[201] = 8'h00;
    mem[202] = 8'hc0;
    mem[203] = 8'h03;
    mem[204] = 8'h80;
    mem[205] = 8'h07;
    mem[206] = 8'h00;
    mem[207] = 8'h00;
    mem[208] = 8'h00;
    mem[209] = 8'h00;
    mem[210] = 8'hc0;
    mem[211] = 8'h03;
    mem[212] = 8'h80;
    mem[213] = 8'h07;
    mem[214] = 8'h00;
    mem[215] = 8'h00;
    mem[216] = 8'h00;
    mem[217] = 8'h00;
    mem[218] = 8'h00;
    mem[219] = 8'h00;
    mem[220] = 8'h80;
    mem[221] = 8'h07;
    mem[222] = 8'h00;
    mem[223] = 8'h00;
    mem[224] = 8'h00;
    mem[225] = 8'h00;
    mem[226] = 8'h00;
    mem[227] = 8'h00;
    mem[228] = 8'h80;
    mem[229] = 8'h07;
    mem[230] = 8'h00;
    mem[231] = 8'h00;
    mem[232] = 8'h00;
    mem[233] = 8'h00;
    mem[234] = 8'h00;
    mem[235] = 8'h00;
    mem[236] = 8'hc0;
    mem[237] = 8'h07;
    mem[238] = 8'h00;
    mem[239] = 8'h00;
    mem[240] = 8'h00;
    mem[241] = 8'h00;
    mem[242] = 8'h00;
    mem[243] = 8'h00;
    mem[244] = 8'hc0;
    mem[245] = 8'h03;
    mem[246] = 8'h00;
    mem[247] = 8'h00;
    mem[248] = 8'h00;
    mem[249] = 8'h00;
    mem[250] = 8'h00;
    mem[251] = 8'h00;
    mem[252] = 8'he0;
    mem[253] = 8'h03;
    mem[254] = 8'h00;
    mem[255] = 8'h00;
    mem[256] = 8'h00;
    mem[257] = 8'h00;
    mem[258] = 8'h00;
    mem[259] = 8'h00;
    mem[260] = 8'hf0;
    mem[261] = 8'h01;
    mem[262] = 8'h00;
    mem[263] = 8'h00;
    mem[264] = 8'h00;
    mem[265] = 8'h00;
    mem[266] = 8'h00;
    mem[267] = 8'h00;
    mem[268] = 8'hf8;
    mem[269] = 8'h00;
    mem[270] = 8'h00;
    mem[271] = 8'h00;
    mem[272] = 8'h00;
    mem[273] = 8'h00;
    mem[274] = 8'h00;
    mem[275] = 8'h00;
    mem[276] = 8'h7c;
    mem[277] = 8'h00;
    mem[278] = 8'h00;
    mem[279] = 8'h00;
    mem[280] = 8'h00;
    mem[281] = 8'h00;
    mem[282] = 8'h00;
    mem[283] = 8'h00;
    mem[284] = 8'h3e;
    mem[285] = 8'h00;
    mem[286] = 8'h00;
    mem[287] = 8'h00;
    mem[288] = 8'h00;
    mem[289] = 8'h00;
    mem[290] = 8'h00;
    mem[291] = 8'h00;
    mem[292] = 8'h3f;
    mem[293] = 8'h00;
    mem[294] = 8'h00;
    mem[295] = 8'h00;
    mem[296] = 8'h00;
    mem[297] = 8'h00;
    mem[298] = 8'h00;
    mem[299] = 8'h80;
    mem[300] = 8'h1f;
    mem[301] = 8'h00;
    mem[302] = 8'h00;
    mem[303] = 8'h00;
    mem[304] = 8'h00;
    mem[305] = 8'h00;
    mem[306] = 8'h00;
    mem[307] = 8'hc0;
    mem[308] = 8'h0f;
    mem[309] = 8'h00;
    mem[310] = 8'h00;
    mem[311] = 8'h00;
    mem[312] = 8'h00;
    mem[313] = 8'h00;
    mem[314] = 8'h00;
    mem[315] = 8'he0;
    mem[316] = 8'h07;
    mem[317] = 8'h00;
    mem[318] = 8'h00;
    mem[319] = 8'h00;
    mem[320] = 8'h00;
    mem[321] = 8'h00;
    mem[322] = 8'h00;
    mem[323] = 8'hf0;
    mem[324] = 8'h03;
    mem[325] = 8'h00;
    mem[326] = 8'h00;
    mem[327] = 8'h00;
    mem[328] = 8'h00;
    mem[329] = 8'h00;
    mem[330] = 8'h00;
    mem[331] = 8'hf8;
    mem[332] = 8'h01;
    mem[333] = 8'h00;
    mem[334] = 8'h00;
    mem[335] = 8'h00;
    mem[336] = 8'h00;
    mem[337] = 8'h00;
    mem[338] = 8'h00;
    mem[339] = 8'hfc;
    mem[340] = 8'h00;
    mem[341] = 8'h00;
    mem[342] = 8'h00;
    mem[343] = 8'h00;
    mem[344] = 8'h00;
    mem[345] = 8'h00;
    mem[346] = 8'h00;
    mem[347] = 8'h3e;
    mem[348] = 8'h00;
    mem[349] = 8'h00;
    mem[350] = 8'h00;
    mem[351] = 8'h00;
    mem[352] = 8'h00;
    mem[353] = 8'h00;
    mem[354] = 8'h00;
    mem[355] = 8'h1f;
    mem[356] = 8'h00;
    mem[357] = 8'h00;
    mem[358] = 8'h00;
    mem[359] = 8'h00;
    mem[360] = 8'h00;
    mem[361] = 8'h00;
    mem[362] = 8'h80;
    mem[363] = 8'h0f;
    mem[364] = 8'h00;
    mem[365] = 8'h00;
    mem[366] = 8'h00;
    mem[367] = 8'h00;
    mem[368] = 8'h00;
    mem[369] = 8'h00;
    mem[370] = 8'hc0;
    mem[371] = 8'h0f;
    mem[372] = 8'h00;
    mem[373] = 8'h00;
    mem[374] = 8'h00;
    mem[375] = 8'h00;
    mem[376] = 8'h00;
    mem[377] = 8'h00;
    mem[378] = 8'he0;
    mem[379] = 8'hff;
    mem[380] = 8'hff;
    mem[381] = 8'h0f;
    mem[382] = 8'h00;
    mem[383] = 8'h00;
    mem[384] = 8'h00;
    mem[385] = 8'h00;
    mem[386] = 8'he0;
    mem[387] = 8'hff;
    mem[388] = 8'hff;
    mem[389] = 8'h0f;
    mem[390] = 8'h00;
    mem[391] = 8'h00;
    mem[392] = 8'h00;
    mem[393] = 8'h00;
    mem[394] = 8'he0;
    mem[395] = 8'hff;
    mem[396] = 8'hff;
    mem[397] = 8'h0f;
    mem[398] = 8'h00;
    mem[399] = 8'h00;
    mem[400] = 8'h00;
    mem[401] = 8'h00;
    mem[402] = 8'h00;
    mem[403] = 8'h00;
    mem[404] = 8'h00;
    mem[405] = 8'h00;
    mem[406] = 8'h00;
    mem[407] = 8'h00;
    mem[408] = 8'h00;
    mem[409] = 8'h00;
    mem[410] = 8'h00;
    mem[411] = 8'h00;
    mem[412] = 8'h00;
    mem[413] = 8'h00;
    mem[414] = 8'h00;
    mem[415] = 8'h00;
    mem[416] = 8'h00;
    mem[417] = 8'h00;
    mem[418] = 8'h00;
    mem[419] = 8'h00;
    mem[420] = 8'h00;
    mem[421] = 8'h00;
    mem[422] = 8'h00;
    mem[423] = 8'h00;
    mem[424] = 8'h00;
    mem[425] = 8'h00;
    mem[426] = 8'h00;
    mem[427] = 8'h00;
    mem[428] = 8'h00;
    mem[429] = 8'h00;
    mem[430] = 8'h00;
    mem[431] = 8'h00;
    mem[432] = 8'h00;
    mem[433] = 8'h00;
    mem[434] = 8'h00;
    mem[435] = 8'h00;
    mem[436] = 8'h00;
    mem[437] = 8'h00;
    mem[438] = 8'h00;
    mem[439] = 8'h00;
    mem[440] = 8'h00;
    mem[441] = 8'h00;
    mem[442] = 8'h00;
    mem[443] = 8'h00;
    mem[444] = 8'h00;
    mem[445] = 8'h00;
    mem[446] = 8'h00;
    mem[447] = 8'h00;
    mem[448] = 8'h00;
    mem[449] = 8'h00;
    mem[450] = 8'h00;
    mem[451] = 8'h00;
    mem[452] = 8'h00;
    mem[453] = 8'h00;
    mem[454] = 8'h00;
    mem[455] = 8'h00;
    mem[456] = 8'h00;
    mem[457] = 8'h00;
    mem[458] = 8'h00;
    mem[459] = 8'h00;
    mem[460] = 8'h00;
    mem[461] = 8'h00;
    mem[462] = 8'h00;
    mem[463] = 8'h00;
    mem[464] = 8'h00;
    mem[465] = 8'h00;
    mem[466] = 8'h00;
    mem[467] = 8'h00;
    mem[468] = 8'h00;
    mem[469] = 8'h00;
    mem[470] = 8'h00;
    mem[471] = 8'h00;
    mem[472] = 8'h00;
    mem[473] = 8'h00;
    mem[474] = 8'h00;
    mem[475] = 8'h00;
    mem[476] = 8'h00;
    mem[477] = 8'h00;
    mem[478] = 8'h00;
    mem[479] = 8'h00;
    mem[480] = 8'h00;
    mem[481] = 8'h00;
    mem[482] = 8'h00;
    mem[483] = 8'h00;
    mem[484] = 8'h00;
    mem[485] = 8'h00;
    mem[486] = 8'h00;
    mem[487] = 8'h00;
    mem[488] = 8'h00;
    mem[489] = 8'h00;
    mem[490] = 8'h00;
    mem[491] = 8'h00;
    mem[492] = 8'h00;
    mem[493] = 8'h00;
    mem[494] = 8'h00;
    mem[495] = 8'h00;
    mem[496] = 8'h00;
    mem[497] = 8'h00;
    mem[498] = 8'h00;
    mem[499] = 8'h00;
    mem[500] = 8'h00;
    mem[501] = 8'h00;
    mem[502] = 8'h00;
    mem[503] = 8'h00;
    mem[504] = 8'h00;
    mem[505] = 8'h00;
    mem[506] = 8'h00;
    mem[507] = 8'h00;
    mem[508] = 8'h00;
    mem[509] = 8'h00;
    mem[510] = 8'h00;
    mem[511] = 8'h00;
  end

  wire [8:0] addr = {y[5:0], x[5:3]};
  assign pixel = mem[addr][x&7];

endmodule

module glyph_4 (
    input wire [5:0] x,
    input wire [5:0] y,
    output wire pixel
);

  reg [7:0] mem[511:0];
  initial begin
    mem[0] = 8'h00;
    mem[1] = 8'h00;
    mem[2] = 8'h00;
    mem[3] = 8'h00;
    mem[4] = 8'h00;
    mem[5] = 8'h00;
    mem[6] = 8'h00;
    mem[7] = 8'h00;
    mem[8] = 8'h00;
    mem[9] = 8'h00;
    mem[10] = 8'h00;
    mem[11] = 8'h00;
    mem[12] = 8'h00;
    mem[13] = 8'h00;
    mem[14] = 8'h00;
    mem[15] = 8'h00;
    mem[16] = 8'h00;
    mem[17] = 8'h00;
    mem[18] = 8'h00;
    mem[19] = 8'h00;
    mem[20] = 8'h00;
    mem[21] = 8'h00;
    mem[22] = 8'h00;
    mem[23] = 8'h00;
    mem[24] = 8'h00;
    mem[25] = 8'h00;
    mem[26] = 8'h00;
    mem[27] = 8'h00;
    mem[28] = 8'h00;
    mem[29] = 8'h00;
    mem[30] = 8'h00;
    mem[31] = 8'h00;
    mem[32] = 8'h00;
    mem[33] = 8'h00;
    mem[34] = 8'h00;
    mem[35] = 8'h00;
    mem[36] = 8'h00;
    mem[37] = 8'h00;
    mem[38] = 8'h00;
    mem[39] = 8'h00;
    mem[40] = 8'h00;
    mem[41] = 8'h00;
    mem[42] = 8'h00;
    mem[43] = 8'h00;
    mem[44] = 8'h00;
    mem[45] = 8'h00;
    mem[46] = 8'h00;
    mem[47] = 8'h00;
    mem[48] = 8'h00;
    mem[49] = 8'h00;
    mem[50] = 8'h00;
    mem[51] = 8'h00;
    mem[52] = 8'h00;
    mem[53] = 8'h00;
    mem[54] = 8'h00;
    mem[55] = 8'h00;
    mem[56] = 8'h00;
    mem[57] = 8'h00;
    mem[58] = 8'h00;
    mem[59] = 8'h00;
    mem[60] = 8'h00;
    mem[61] = 8'h00;
    mem[62] = 8'h00;
    mem[63] = 8'h00;
    mem[64] = 8'h00;
    mem[65] = 8'h00;
    mem[66] = 8'h00;
    mem[67] = 8'h00;
    mem[68] = 8'h00;
    mem[69] = 8'h00;
    mem[70] = 8'h00;
    mem[71] = 8'h00;
    mem[72] = 8'h00;
    mem[73] = 8'h00;
    mem[74] = 8'h00;
    mem[75] = 8'h00;
    mem[76] = 8'h00;
    mem[77] = 8'h00;
    mem[78] = 8'h00;
    mem[79] = 8'h00;
    mem[80] = 8'h00;
    mem[81] = 8'h00;
    mem[82] = 8'h00;
    mem[83] = 8'h00;
    mem[84] = 8'h00;
    mem[85] = 8'h00;
    mem[86] = 8'h00;
    mem[87] = 8'h00;
    mem[88] = 8'h00;
    mem[89] = 8'h00;
    mem[90] = 8'h00;
    mem[91] = 8'h00;
    mem[92] = 8'h00;
    mem[93] = 8'h00;
    mem[94] = 8'h00;
    mem[95] = 8'h00;
    mem[96] = 8'h00;
    mem[97] = 8'h00;
    mem[98] = 8'h00;
    mem[99] = 8'h00;
    mem[100] = 8'h00;
    mem[101] = 8'h00;
    mem[102] = 8'h00;
    mem[103] = 8'h00;
    mem[104] = 8'h00;
    mem[105] = 8'h00;
    mem[106] = 8'h00;
    mem[107] = 8'h00;
    mem[108] = 8'h00;
    mem[109] = 8'h00;
    mem[110] = 8'h00;
    mem[111] = 8'h00;
    mem[112] = 8'h00;
    mem[113] = 8'h00;
    mem[114] = 8'h00;
    mem[115] = 8'h00;
    mem[116] = 8'h00;
    mem[117] = 8'h00;
    mem[118] = 8'h00;
    mem[119] = 8'h00;
    mem[120] = 8'h00;
    mem[121] = 8'h00;
    mem[122] = 8'h00;
    mem[123] = 8'h00;
    mem[124] = 8'h00;
    mem[125] = 8'h00;
    mem[126] = 8'h00;
    mem[127] = 8'h00;
    mem[128] = 8'h00;
    mem[129] = 8'h00;
    mem[130] = 8'h00;
    mem[131] = 8'h00;
    mem[132] = 8'h00;
    mem[133] = 8'h00;
    mem[134] = 8'h00;
    mem[135] = 8'h00;
    mem[136] = 8'h00;
    mem[137] = 8'h00;
    mem[138] = 8'h00;
    mem[139] = 8'h00;
    mem[140] = 8'hf0;
    mem[141] = 8'h01;
    mem[142] = 8'h00;
    mem[143] = 8'h00;
    mem[144] = 8'h00;
    mem[145] = 8'h00;
    mem[146] = 8'h00;
    mem[147] = 8'h00;
    mem[148] = 8'hf8;
    mem[149] = 8'h01;
    mem[150] = 8'h00;
    mem[151] = 8'h00;
    mem[152] = 8'h00;
    mem[153] = 8'h00;
    mem[154] = 8'h00;
    mem[155] = 8'h00;
    mem[156] = 8'hfc;
    mem[157] = 8'h01;
    mem[158] = 8'h00;
    mem[159] = 8'h00;
    mem[160] = 8'h00;
    mem[161] = 8'h00;
    mem[162] = 8'h00;
    mem[163] = 8'h00;
    mem[164] = 8'hfc;
    mem[165] = 8'h01;
    mem[166] = 8'h00;
    mem[167] = 8'h00;
    mem[168] = 8'h00;
    mem[169] = 8'h00;
    mem[170] = 8'h00;
    mem[171] = 8'h00;
    mem[172] = 8'hfe;
    mem[173] = 8'h01;
    mem[174] = 8'h00;
    mem[175] = 8'h00;
    mem[176] = 8'h00;
    mem[177] = 8'h00;
    mem[178] = 8'h00;
    mem[179] = 8'h00;
    mem[180] = 8'hff;
    mem[181] = 8'h01;
    mem[182] = 8'h00;
    mem[183] = 8'h00;
    mem[184] = 8'h00;
    mem[185] = 8'h00;
    mem[186] = 8'h00;
    mem[187] = 8'h80;
    mem[188] = 8'hf7;
    mem[189] = 8'h01;
    mem[190] = 8'h00;
    mem[191] = 8'h00;
    mem[192] = 8'h00;
    mem[193] = 8'h00;
    mem[194] = 8'h00;
    mem[195] = 8'h80;
    mem[196] = 8'hf7;
    mem[197] = 8'h01;
    mem[198] = 8'h00;
    mem[199] = 8'h00;
    mem[200] = 8'h00;
    mem[201] = 8'h00;
    mem[202] = 8'h00;
    mem[203] = 8'hc0;
    mem[204] = 8'hf3;
    mem[205] = 8'h01;
    mem[206] = 8'h00;
    mem[207] = 8'h00;
    mem[208] = 8'h00;
    mem[209] = 8'h00;
    mem[210] = 8'h00;
    mem[211] = 8'he0;
    mem[212] = 8'hf3;
    mem[213] = 8'h01;
    mem[214] = 8'h00;
    mem[215] = 8'h00;
    mem[216] = 8'h00;
    mem[217] = 8'h00;
    mem[218] = 8'h00;
    mem[219] = 8'he0;
    mem[220] = 8'hf1;
    mem[221] = 8'h01;
    mem[222] = 8'h00;
    mem[223] = 8'h00;
    mem[224] = 8'h00;
    mem[225] = 8'h00;
    mem[226] = 8'h00;
    mem[227] = 8'hf0;
    mem[228] = 8'hf0;
    mem[229] = 8'h01;
    mem[230] = 8'h00;
    mem[231] = 8'h00;
    mem[232] = 8'h00;
    mem[233] = 8'h00;
    mem[234] = 8'h00;
    mem[235] = 8'hf8;
    mem[236] = 8'hf0;
    mem[237] = 8'h01;
    mem[238] = 8'h00;
    mem[239] = 8'h00;
    mem[240] = 8'h00;
    mem[241] = 8'h00;
    mem[242] = 8'h00;
    mem[243] = 8'h78;
    mem[244] = 8'hf0;
    mem[245] = 8'h01;
    mem[246] = 8'h00;
    mem[247] = 8'h00;
    mem[248] = 8'h00;
    mem[249] = 8'h00;
    mem[250] = 8'h00;
    mem[251] = 8'h3c;
    mem[252] = 8'hf0;
    mem[253] = 8'h01;
    mem[254] = 8'h00;
    mem[255] = 8'h00;
    mem[256] = 8'h00;
    mem[257] = 8'h00;
    mem[258] = 8'h00;
    mem[259] = 8'h1e;
    mem[260] = 8'hf0;
    mem[261] = 8'h01;
    mem[262] = 8'h00;
    mem[263] = 8'h00;
    mem[264] = 8'h00;
    mem[265] = 8'h00;
    mem[266] = 8'h00;
    mem[267] = 8'h1e;
    mem[268] = 8'hf0;
    mem[269] = 8'h01;
    mem[270] = 8'h00;
    mem[271] = 8'h00;
    mem[272] = 8'h00;
    mem[273] = 8'h00;
    mem[274] = 8'h00;
    mem[275] = 8'h0f;
    mem[276] = 8'hf0;
    mem[277] = 8'h01;
    mem[278] = 8'h00;
    mem[279] = 8'h00;
    mem[280] = 8'h00;
    mem[281] = 8'h00;
    mem[282] = 8'h80;
    mem[283] = 8'h07;
    mem[284] = 8'hf0;
    mem[285] = 8'h01;
    mem[286] = 8'h00;
    mem[287] = 8'h00;
    mem[288] = 8'h00;
    mem[289] = 8'h00;
    mem[290] = 8'hc0;
    mem[291] = 8'h07;
    mem[292] = 8'hf0;
    mem[293] = 8'h01;
    mem[294] = 8'h00;
    mem[295] = 8'h00;
    mem[296] = 8'h00;
    mem[297] = 8'h00;
    mem[298] = 8'hc0;
    mem[299] = 8'h03;
    mem[300] = 8'hf0;
    mem[301] = 8'h01;
    mem[302] = 8'h00;
    mem[303] = 8'h00;
    mem[304] = 8'h00;
    mem[305] = 8'h00;
    mem[306] = 8'he0;
    mem[307] = 8'h01;
    mem[308] = 8'hf0;
    mem[309] = 8'h01;
    mem[310] = 8'h00;
    mem[311] = 8'h00;
    mem[312] = 8'h00;
    mem[313] = 8'h00;
    mem[314] = 8'hf0;
    mem[315] = 8'hff;
    mem[316] = 8'hff;
    mem[317] = 8'h1f;
    mem[318] = 8'h00;
    mem[319] = 8'h00;
    mem[320] = 8'h00;
    mem[321] = 8'h00;
    mem[322] = 8'hf0;
    mem[323] = 8'hff;
    mem[324] = 8'hff;
    mem[325] = 8'h1f;
    mem[326] = 8'h00;
    mem[327] = 8'h00;
    mem[328] = 8'h00;
    mem[329] = 8'h00;
    mem[330] = 8'hf0;
    mem[331] = 8'hff;
    mem[332] = 8'hff;
    mem[333] = 8'h1f;
    mem[334] = 8'h00;
    mem[335] = 8'h00;
    mem[336] = 8'h00;
    mem[337] = 8'h00;
    mem[338] = 8'h00;
    mem[339] = 8'h00;
    mem[340] = 8'hf0;
    mem[341] = 8'h01;
    mem[342] = 8'h00;
    mem[343] = 8'h00;
    mem[344] = 8'h00;
    mem[345] = 8'h00;
    mem[346] = 8'h00;
    mem[347] = 8'h00;
    mem[348] = 8'hf0;
    mem[349] = 8'h01;
    mem[350] = 8'h00;
    mem[351] = 8'h00;
    mem[352] = 8'h00;
    mem[353] = 8'h00;
    mem[354] = 8'h00;
    mem[355] = 8'h00;
    mem[356] = 8'hf0;
    mem[357] = 8'h01;
    mem[358] = 8'h00;
    mem[359] = 8'h00;
    mem[360] = 8'h00;
    mem[361] = 8'h00;
    mem[362] = 8'h00;
    mem[363] = 8'h00;
    mem[364] = 8'hf0;
    mem[365] = 8'h01;
    mem[366] = 8'h00;
    mem[367] = 8'h00;
    mem[368] = 8'h00;
    mem[369] = 8'h00;
    mem[370] = 8'h00;
    mem[371] = 8'h00;
    mem[372] = 8'hf0;
    mem[373] = 8'h01;
    mem[374] = 8'h00;
    mem[375] = 8'h00;
    mem[376] = 8'h00;
    mem[377] = 8'h00;
    mem[378] = 8'h00;
    mem[379] = 8'h00;
    mem[380] = 8'hf0;
    mem[381] = 8'h01;
    mem[382] = 8'h00;
    mem[383] = 8'h00;
    mem[384] = 8'h00;
    mem[385] = 8'h00;
    mem[386] = 8'h00;
    mem[387] = 8'h00;
    mem[388] = 8'hf0;
    mem[389] = 8'h01;
    mem[390] = 8'h00;
    mem[391] = 8'h00;
    mem[392] = 8'h00;
    mem[393] = 8'h00;
    mem[394] = 8'h00;
    mem[395] = 8'h00;
    mem[396] = 8'hf0;
    mem[397] = 8'h01;
    mem[398] = 8'h00;
    mem[399] = 8'h00;
    mem[400] = 8'h00;
    mem[401] = 8'h00;
    mem[402] = 8'h00;
    mem[403] = 8'h00;
    mem[404] = 8'h00;
    mem[405] = 8'h00;
    mem[406] = 8'h00;
    mem[407] = 8'h00;
    mem[408] = 8'h00;
    mem[409] = 8'h00;
    mem[410] = 8'h00;
    mem[411] = 8'h00;
    mem[412] = 8'h00;
    mem[413] = 8'h00;
    mem[414] = 8'h00;
    mem[415] = 8'h00;
    mem[416] = 8'h00;
    mem[417] = 8'h00;
    mem[418] = 8'h00;
    mem[419] = 8'h00;
    mem[420] = 8'h00;
    mem[421] = 8'h00;
    mem[422] = 8'h00;
    mem[423] = 8'h00;
    mem[424] = 8'h00;
    mem[425] = 8'h00;
    mem[426] = 8'h00;
    mem[427] = 8'h00;
    mem[428] = 8'h00;
    mem[429] = 8'h00;
    mem[430] = 8'h00;
    mem[431] = 8'h00;
    mem[432] = 8'h00;
    mem[433] = 8'h00;
    mem[434] = 8'h00;
    mem[435] = 8'h00;
    mem[436] = 8'h00;
    mem[437] = 8'h00;
    mem[438] = 8'h00;
    mem[439] = 8'h00;
    mem[440] = 8'h00;
    mem[441] = 8'h00;
    mem[442] = 8'h00;
    mem[443] = 8'h00;
    mem[444] = 8'h00;
    mem[445] = 8'h00;
    mem[446] = 8'h00;
    mem[447] = 8'h00;
    mem[448] = 8'h00;
    mem[449] = 8'h00;
    mem[450] = 8'h00;
    mem[451] = 8'h00;
    mem[452] = 8'h00;
    mem[453] = 8'h00;
    mem[454] = 8'h00;
    mem[455] = 8'h00;
    mem[456] = 8'h00;
    mem[457] = 8'h00;
    mem[458] = 8'h00;
    mem[459] = 8'h00;
    mem[460] = 8'h00;
    mem[461] = 8'h00;
    mem[462] = 8'h00;
    mem[463] = 8'h00;
    mem[464] = 8'h00;
    mem[465] = 8'h00;
    mem[466] = 8'h00;
    mem[467] = 8'h00;
    mem[468] = 8'h00;
    mem[469] = 8'h00;
    mem[470] = 8'h00;
    mem[471] = 8'h00;
    mem[472] = 8'h00;
    mem[473] = 8'h00;
    mem[474] = 8'h00;
    mem[475] = 8'h00;
    mem[476] = 8'h00;
    mem[477] = 8'h00;
    mem[478] = 8'h00;
    mem[479] = 8'h00;
    mem[480] = 8'h00;
    mem[481] = 8'h00;
    mem[482] = 8'h00;
    mem[483] = 8'h00;
    mem[484] = 8'h00;
    mem[485] = 8'h00;
    mem[486] = 8'h00;
    mem[487] = 8'h00;
    mem[488] = 8'h00;
    mem[489] = 8'h00;
    mem[490] = 8'h00;
    mem[491] = 8'h00;
    mem[492] = 8'h00;
    mem[493] = 8'h00;
    mem[494] = 8'h00;
    mem[495] = 8'h00;
    mem[496] = 8'h00;
    mem[497] = 8'h00;
    mem[498] = 8'h00;
    mem[499] = 8'h00;
    mem[500] = 8'h00;
    mem[501] = 8'h00;
    mem[502] = 8'h00;
    mem[503] = 8'h00;
    mem[504] = 8'h00;
    mem[505] = 8'h00;
    mem[506] = 8'h00;
    mem[507] = 8'h00;
    mem[508] = 8'h00;
    mem[509] = 8'h00;
    mem[510] = 8'h00;
    mem[511] = 8'h00;
  end

  wire [8:0] addr = {y[5:0], x[5:3]};
  assign pixel = mem[addr][x&7];

endmodule

module glyph_8 (
    input wire [5:0] x,
    input wire [5:0] y,
    output wire pixel
);

  reg [7:0] mem[511:0];
  initial begin
    mem[0] = 8'h00;
    mem[1] = 8'h00;
    mem[2] = 8'h00;
    mem[3] = 8'h00;
    mem[4] = 8'h00;
    mem[5] = 8'h00;
    mem[6] = 8'h00;
    mem[7] = 8'h00;
    mem[8] = 8'h00;
    mem[9] = 8'h00;
    mem[10] = 8'h00;
    mem[11] = 8'h00;
    mem[12] = 8'h00;
    mem[13] = 8'h00;
    mem[14] = 8'h00;
    mem[15] = 8'h00;
    mem[16] = 8'h00;
    mem[17] = 8'h00;
    mem[18] = 8'h00;
    mem[19] = 8'h00;
    mem[20] = 8'h00;
    mem[21] = 8'h00;
    mem[22] = 8'h00;
    mem[23] = 8'h00;
    mem[24] = 8'h00;
    mem[25] = 8'h00;
    mem[26] = 8'h00;
    mem[27] = 8'h00;
    mem[28] = 8'h00;
    mem[29] = 8'h00;
    mem[30] = 8'h00;
    mem[31] = 8'h00;
    mem[32] = 8'h00;
    mem[33] = 8'h00;
    mem[34] = 8'h00;
    mem[35] = 8'h00;
    mem[36] = 8'h00;
    mem[37] = 8'h00;
    mem[38] = 8'h00;
    mem[39] = 8'h00;
    mem[40] = 8'h00;
    mem[41] = 8'h00;
    mem[42] = 8'h00;
    mem[43] = 8'h00;
    mem[44] = 8'h00;
    mem[45] = 8'h00;
    mem[46] = 8'h00;
    mem[47] = 8'h00;
    mem[48] = 8'h00;
    mem[49] = 8'h00;
    mem[50] = 8'h00;
    mem[51] = 8'h00;
    mem[52] = 8'h00;
    mem[53] = 8'h00;
    mem[54] = 8'h00;
    mem[55] = 8'h00;
    mem[56] = 8'h00;
    mem[57] = 8'h00;
    mem[58] = 8'h00;
    mem[59] = 8'h00;
    mem[60] = 8'h00;
    mem[61] = 8'h00;
    mem[62] = 8'h00;
    mem[63] = 8'h00;
    mem[64] = 8'h00;
    mem[65] = 8'h00;
    mem[66] = 8'h00;
    mem[67] = 8'h00;
    mem[68] = 8'h00;
    mem[69] = 8'h00;
    mem[70] = 8'h00;
    mem[71] = 8'h00;
    mem[72] = 8'h00;
    mem[73] = 8'h00;
    mem[74] = 8'h00;
    mem[75] = 8'h00;
    mem[76] = 8'h00;
    mem[77] = 8'h00;
    mem[78] = 8'h00;
    mem[79] = 8'h00;
    mem[80] = 8'h00;
    mem[81] = 8'h00;
    mem[82] = 8'h00;
    mem[83] = 8'h00;
    mem[84] = 8'h00;
    mem[85] = 8'h00;
    mem[86] = 8'h00;
    mem[87] = 8'h00;
    mem[88] = 8'h00;
    mem[89] = 8'h00;
    mem[90] = 8'h00;
    mem[91] = 8'h00;
    mem[92] = 8'h00;
    mem[93] = 8'h00;
    mem[94] = 8'h00;
    mem[95] = 8'h00;
    mem[96] = 8'h00;
    mem[97] = 8'h00;
    mem[98] = 8'h00;
    mem[99] = 8'h00;
    mem[100] = 8'h00;
    mem[101] = 8'h00;
    mem[102] = 8'h00;
    mem[103] = 8'h00;
    mem[104] = 8'h00;
    mem[105] = 8'h00;
    mem[106] = 8'h00;
    mem[107] = 8'h00;
    mem[108] = 8'h00;
    mem[109] = 8'h00;
    mem[110] = 8'h00;
    mem[111] = 8'h00;
    mem[112] = 8'h00;
    mem[113] = 8'h00;
    mem[114] = 8'h00;
    mem[115] = 8'h00;
    mem[116] = 8'h00;
    mem[117] = 8'h00;
    mem[118] = 8'h00;
    mem[119] = 8'h00;
    mem[120] = 8'h00;
    mem[121] = 8'h00;
    mem[122] = 8'h00;
    mem[123] = 8'h00;
    mem[124] = 8'h00;
    mem[125] = 8'h00;
    mem[126] = 8'h00;
    mem[127] = 8'h00;
    mem[128] = 8'h00;
    mem[129] = 8'h00;
    mem[130] = 8'h00;
    mem[131] = 8'h00;
    mem[132] = 8'h00;
    mem[133] = 8'h00;
    mem[134] = 8'h00;
    mem[135] = 8'h00;
    mem[136] = 8'h00;
    mem[137] = 8'h00;
    mem[138] = 8'h00;
    mem[139] = 8'hf8;
    mem[140] = 8'h3f;
    mem[141] = 8'h00;
    mem[142] = 8'h00;
    mem[143] = 8'h00;
    mem[144] = 8'h00;
    mem[145] = 8'h00;
    mem[146] = 8'h00;
    mem[147] = 8'hfe;
    mem[148] = 8'h7f;
    mem[149] = 8'h00;
    mem[150] = 8'h00;
    mem[151] = 8'h00;
    mem[152] = 8'h00;
    mem[153] = 8'h00;
    mem[154] = 8'h00;
    mem[155] = 8'hff;
    mem[156] = 8'hff;
    mem[157] = 8'h01;
    mem[158] = 8'h00;
    mem[159] = 8'h00;
    mem[160] = 8'h00;
    mem[161] = 8'h00;
    mem[162] = 8'h80;
    mem[163] = 8'h1f;
    mem[164] = 8'hf0;
    mem[165] = 8'h03;
    mem[166] = 8'h00;
    mem[167] = 8'h00;
    mem[168] = 8'h00;
    mem[169] = 8'h00;
    mem[170] = 8'hc0;
    mem[171] = 8'h07;
    mem[172] = 8'he0;
    mem[173] = 8'h03;
    mem[174] = 8'h00;
    mem[175] = 8'h00;
    mem[176] = 8'h00;
    mem[177] = 8'h00;
    mem[178] = 8'hc0;
    mem[179] = 8'h07;
    mem[180] = 8'hc0;
    mem[181] = 8'h07;
    mem[182] = 8'h00;
    mem[183] = 8'h00;
    mem[184] = 8'h00;
    mem[185] = 8'h00;
    mem[186] = 8'hc0;
    mem[187] = 8'h03;
    mem[188] = 8'hc0;
    mem[189] = 8'h07;
    mem[190] = 8'h00;
    mem[191] = 8'h00;
    mem[192] = 8'h00;
    mem[193] = 8'h00;
    mem[194] = 8'hc0;
    mem[195] = 8'h03;
    mem[196] = 8'hc0;
    mem[197] = 8'h07;
    mem[198] = 8'h00;
    mem[199] = 8'h00;
    mem[200] = 8'h00;
    mem[201] = 8'h00;
    mem[202] = 8'hc0;
    mem[203] = 8'h03;
    mem[204] = 8'hc0;
    mem[205] = 8'h07;
    mem[206] = 8'h00;
    mem[207] = 8'h00;
    mem[208] = 8'h00;
    mem[209] = 8'h00;
    mem[210] = 8'hc0;
    mem[211] = 8'h03;
    mem[212] = 8'hc0;
    mem[213] = 8'h07;
    mem[214] = 8'h00;
    mem[215] = 8'h00;
    mem[216] = 8'h00;
    mem[217] = 8'h00;
    mem[218] = 8'hc0;
    mem[219] = 8'h03;
    mem[220] = 8'hc0;
    mem[221] = 8'h07;
    mem[222] = 8'h00;
    mem[223] = 8'h00;
    mem[224] = 8'h00;
    mem[225] = 8'h00;
    mem[226] = 8'hc0;
    mem[227] = 8'h07;
    mem[228] = 8'hc0;
    mem[229] = 8'h03;
    mem[230] = 8'h00;
    mem[231] = 8'h00;
    mem[232] = 8'h00;
    mem[233] = 8'h00;
    mem[234] = 8'h80;
    mem[235] = 8'h0f;
    mem[236] = 8'he0;
    mem[237] = 8'h03;
    mem[238] = 8'h00;
    mem[239] = 8'h00;
    mem[240] = 8'h00;
    mem[241] = 8'h00;
    mem[242] = 8'h00;
    mem[243] = 8'h1f;
    mem[244] = 8'hf8;
    mem[245] = 8'h01;
    mem[246] = 8'h00;
    mem[247] = 8'h00;
    mem[248] = 8'h00;
    mem[249] = 8'h00;
    mem[250] = 8'h00;
    mem[251] = 8'hfe;
    mem[252] = 8'hff;
    mem[253] = 8'h00;
    mem[254] = 8'h00;
    mem[255] = 8'h00;
    mem[256] = 8'h00;
    mem[257] = 8'h00;
    mem[258] = 8'h00;
    mem[259] = 8'hfc;
    mem[260] = 8'h3f;
    mem[261] = 8'h00;
    mem[262] = 8'h00;
    mem[263] = 8'h00;
    mem[264] = 8'h00;
    mem[265] = 8'h00;
    mem[266] = 8'h00;
    mem[267] = 8'hff;
    mem[268] = 8'hff;
    mem[269] = 8'h00;
    mem[270] = 8'h00;
    mem[271] = 8'h00;
    mem[272] = 8'h00;
    mem[273] = 8'h00;
    mem[274] = 8'h80;
    mem[275] = 8'h1f;
    mem[276] = 8'hfc;
    mem[277] = 8'h01;
    mem[278] = 8'h00;
    mem[279] = 8'h00;
    mem[280] = 8'h00;
    mem[281] = 8'h00;
    mem[282] = 8'hc0;
    mem[283] = 8'h07;
    mem[284] = 8'he0;
    mem[285] = 8'h03;
    mem[286] = 8'h00;
    mem[287] = 8'h00;
    mem[288] = 8'h00;
    mem[289] = 8'h00;
    mem[290] = 8'he0;
    mem[291] = 8'h03;
    mem[292] = 8'hc0;
    mem[293] = 8'h03;
    mem[294] = 8'h00;
    mem[295] = 8'h00;
    mem[296] = 8'h00;
    mem[297] = 8'h00;
    mem[298] = 8'he0;
    mem[299] = 8'h01;
    mem[300] = 8'hc0;
    mem[301] = 8'h07;
    mem[302] = 8'h00;
    mem[303] = 8'h00;
    mem[304] = 8'h00;
    mem[305] = 8'h00;
    mem[306] = 8'hf0;
    mem[307] = 8'h01;
    mem[308] = 8'h80;
    mem[309] = 8'h07;
    mem[310] = 8'h00;
    mem[311] = 8'h00;
    mem[312] = 8'h00;
    mem[313] = 8'h00;
    mem[314] = 8'hf0;
    mem[315] = 8'h01;
    mem[316] = 8'h80;
    mem[317] = 8'h07;
    mem[318] = 8'h00;
    mem[319] = 8'h00;
    mem[320] = 8'h00;
    mem[321] = 8'h00;
    mem[322] = 8'hf0;
    mem[323] = 8'h01;
    mem[324] = 8'h80;
    mem[325] = 8'h07;
    mem[326] = 8'h00;
    mem[327] = 8'h00;
    mem[328] = 8'h00;
    mem[329] = 8'h00;
    mem[330] = 8'hf0;
    mem[331] = 8'h01;
    mem[332] = 8'h80;
    mem[333] = 8'h07;
    mem[334] = 8'h00;
    mem[335] = 8'h00;
    mem[336] = 8'h00;
    mem[337] = 8'h00;
    mem[338] = 8'hf0;
    mem[339] = 8'h01;
    mem[340] = 8'h80;
    mem[341] = 8'h07;
    mem[342] = 8'h00;
    mem[343] = 8'h00;
    mem[344] = 8'h00;
    mem[345] = 8'h00;
    mem[346] = 8'hf0;
    mem[347] = 8'h01;
    mem[348] = 8'hc0;
    mem[349] = 8'h07;
    mem[350] = 8'h00;
    mem[351] = 8'h00;
    mem[352] = 8'h00;
    mem[353] = 8'h00;
    mem[354] = 8'he0;
    mem[355] = 8'h03;
    mem[356] = 8'hc0;
    mem[357] = 8'h07;
    mem[358] = 8'h00;
    mem[359] = 8'h00;
    mem[360] = 8'h00;
    mem[361] = 8'h00;
    mem[362] = 8'he0;
    mem[363] = 8'h03;
    mem[364] = 8'he0;
    mem[365] = 8'h03;
    mem[366] = 8'h00;
    mem[367] = 8'h00;
    mem[368] = 8'h00;
    mem[369] = 8'h00;
    mem[370] = 8'hc0;
    mem[371] = 8'h0f;
    mem[372] = 8'hf0;
    mem[373] = 8'h03;
    mem[374] = 8'h00;
    mem[375] = 8'h00;
    mem[376] = 8'h00;
    mem[377] = 8'h00;
    mem[378] = 8'h80;
    mem[379] = 8'hff;
    mem[380] = 8'hff;
    mem[381] = 8'h01;
    mem[382] = 8'h00;
    mem[383] = 8'h00;
    mem[384] = 8'h00;
    mem[385] = 8'h00;
    mem[386] = 8'h00;
    mem[387] = 8'hff;
    mem[388] = 8'h7f;
    mem[389] = 8'h00;
    mem[390] = 8'h00;
    mem[391] = 8'h00;
    mem[392] = 8'h00;
    mem[393] = 8'h00;
    mem[394] = 8'h00;
    mem[395] = 8'hfc;
    mem[396] = 8'h1f;
    mem[397] = 8'h00;
    mem[398] = 8'h00;
    mem[399] = 8'h00;
    mem[400] = 8'h00;
    mem[401] = 8'h00;
    mem[402] = 8'h00;
    mem[403] = 8'h00;
    mem[404] = 8'h00;
    mem[405] = 8'h00;
    mem[406] = 8'h00;
    mem[407] = 8'h00;
    mem[408] = 8'h00;
    mem[409] = 8'h00;
    mem[410] = 8'h00;
    mem[411] = 8'h00;
    mem[412] = 8'h00;
    mem[413] = 8'h00;
    mem[414] = 8'h00;
    mem[415] = 8'h00;
    mem[416] = 8'h00;
    mem[417] = 8'h00;
    mem[418] = 8'h00;
    mem[419] = 8'h00;
    mem[420] = 8'h00;
    mem[421] = 8'h00;
    mem[422] = 8'h00;
    mem[423] = 8'h00;
    mem[424] = 8'h00;
    mem[425] = 8'h00;
    mem[426] = 8'h00;
    mem[427] = 8'h00;
    mem[428] = 8'h00;
    mem[429] = 8'h00;
    mem[430] = 8'h00;
    mem[431] = 8'h00;
    mem[432] = 8'h00;
    mem[433] = 8'h00;
    mem[434] = 8'h00;
    mem[435] = 8'h00;
    mem[436] = 8'h00;
    mem[437] = 8'h00;
    mem[438] = 8'h00;
    mem[439] = 8'h00;
    mem[440] = 8'h00;
    mem[441] = 8'h00;
    mem[442] = 8'h00;
    mem[443] = 8'h00;
    mem[444] = 8'h00;
    mem[445] = 8'h00;
    mem[446] = 8'h00;
    mem[447] = 8'h00;
    mem[448] = 8'h00;
    mem[449] = 8'h00;
    mem[450] = 8'h00;
    mem[451] = 8'h00;
    mem[452] = 8'h00;
    mem[453] = 8'h00;
    mem[454] = 8'h00;
    mem[455] = 8'h00;
    mem[456] = 8'h00;
    mem[457] = 8'h00;
    mem[458] = 8'h00;
    mem[459] = 8'h00;
    mem[460] = 8'h00;
    mem[461] = 8'h00;
    mem[462] = 8'h00;
    mem[463] = 8'h00;
    mem[464] = 8'h00;
    mem[465] = 8'h00;
    mem[466] = 8'h00;
    mem[467] = 8'h00;
    mem[468] = 8'h00;
    mem[469] = 8'h00;
    mem[470] = 8'h00;
    mem[471] = 8'h00;
    mem[472] = 8'h00;
    mem[473] = 8'h00;
    mem[474] = 8'h00;
    mem[475] = 8'h00;
    mem[476] = 8'h00;
    mem[477] = 8'h00;
    mem[478] = 8'h00;
    mem[479] = 8'h00;
    mem[480] = 8'h00;
    mem[481] = 8'h00;
    mem[482] = 8'h00;
    mem[483] = 8'h00;
    mem[484] = 8'h00;
    mem[485] = 8'h00;
    mem[486] = 8'h00;
    mem[487] = 8'h00;
    mem[488] = 8'h00;
    mem[489] = 8'h00;
    mem[490] = 8'h00;
    mem[491] = 8'h00;
    mem[492] = 8'h00;
    mem[493] = 8'h00;
    mem[494] = 8'h00;
    mem[495] = 8'h00;
    mem[496] = 8'h00;
    mem[497] = 8'h00;
    mem[498] = 8'h00;
    mem[499] = 8'h00;
    mem[500] = 8'h00;
    mem[501] = 8'h00;
    mem[502] = 8'h00;
    mem[503] = 8'h00;
    mem[504] = 8'h00;
    mem[505] = 8'h00;
    mem[506] = 8'h00;
    mem[507] = 8'h00;
    mem[508] = 8'h00;
    mem[509] = 8'h00;
    mem[510] = 8'h00;
    mem[511] = 8'h00;
  end

  wire [8:0] addr = {y[5:0], x[5:3]};
  assign pixel = mem[addr][x&7];

endmodule

module glyph_16 (
    input wire [5:0] x,
    input wire [5:0] y,
    output wire pixel
);

  reg [7:0] mem[511:0];
  initial begin
    mem[0] = 8'h00;
    mem[1] = 8'h00;
    mem[2] = 8'h00;
    mem[3] = 8'h00;
    mem[4] = 8'h00;
    mem[5] = 8'h00;
    mem[6] = 8'h00;
    mem[7] = 8'h00;
    mem[8] = 8'h00;
    mem[9] = 8'h00;
    mem[10] = 8'h00;
    mem[11] = 8'h00;
    mem[12] = 8'h00;
    mem[13] = 8'h00;
    mem[14] = 8'h00;
    mem[15] = 8'h00;
    mem[16] = 8'h00;
    mem[17] = 8'h00;
    mem[18] = 8'h00;
    mem[19] = 8'h00;
    mem[20] = 8'h00;
    mem[21] = 8'h00;
    mem[22] = 8'h00;
    mem[23] = 8'h00;
    mem[24] = 8'h00;
    mem[25] = 8'h00;
    mem[26] = 8'h00;
    mem[27] = 8'h00;
    mem[28] = 8'h00;
    mem[29] = 8'h00;
    mem[30] = 8'h00;
    mem[31] = 8'h00;
    mem[32] = 8'h00;
    mem[33] = 8'h00;
    mem[34] = 8'h00;
    mem[35] = 8'h00;
    mem[36] = 8'h00;
    mem[37] = 8'h00;
    mem[38] = 8'h00;
    mem[39] = 8'h00;
    mem[40] = 8'h00;
    mem[41] = 8'h00;
    mem[42] = 8'h00;
    mem[43] = 8'h00;
    mem[44] = 8'h00;
    mem[45] = 8'h00;
    mem[46] = 8'h00;
    mem[47] = 8'h00;
    mem[48] = 8'h00;
    mem[49] = 8'h00;
    mem[50] = 8'h00;
    mem[51] = 8'h00;
    mem[52] = 8'h00;
    mem[53] = 8'h00;
    mem[54] = 8'h00;
    mem[55] = 8'h00;
    mem[56] = 8'h00;
    mem[57] = 8'h00;
    mem[58] = 8'h00;
    mem[59] = 8'h00;
    mem[60] = 8'h00;
    mem[61] = 8'h00;
    mem[62] = 8'h00;
    mem[63] = 8'h00;
    mem[64] = 8'h00;
    mem[65] = 8'h00;
    mem[66] = 8'h00;
    mem[67] = 8'h00;
    mem[68] = 8'h00;
    mem[69] = 8'h00;
    mem[70] = 8'h00;
    mem[71] = 8'h00;
    mem[72] = 8'h00;
    mem[73] = 8'h00;
    mem[74] = 8'h00;
    mem[75] = 8'h00;
    mem[76] = 8'h00;
    mem[77] = 8'h00;
    mem[78] = 8'h00;
    mem[79] = 8'h00;
    mem[80] = 8'h00;
    mem[81] = 8'h00;
    mem[82] = 8'h00;
    mem[83] = 8'h00;
    mem[84] = 8'h00;
    mem[85] = 8'h00;
    mem[86] = 8'h00;
    mem[87] = 8'h00;
    mem[88] = 8'h00;
    mem[89] = 8'h00;
    mem[90] = 8'h00;
    mem[91] = 8'h00;
    mem[92] = 8'h00;
    mem[93] = 8'h00;
    mem[94] = 8'h00;
    mem[95] = 8'h00;
    mem[96] = 8'h00;
    mem[97] = 8'h00;
    mem[98] = 8'h00;
    mem[99] = 8'h00;
    mem[100] = 8'h00;
    mem[101] = 8'h00;
    mem[102] = 8'h00;
    mem[103] = 8'h00;
    mem[104] = 8'h00;
    mem[105] = 8'h00;
    mem[106] = 8'h00;
    mem[107] = 8'h00;
    mem[108] = 8'h00;
    mem[109] = 8'h00;
    mem[110] = 8'h00;
    mem[111] = 8'h00;
    mem[112] = 8'h00;
    mem[113] = 8'h00;
    mem[114] = 8'h00;
    mem[115] = 8'h00;
    mem[116] = 8'h00;
    mem[117] = 8'h00;
    mem[118] = 8'h00;
    mem[119] = 8'h00;
    mem[120] = 8'h00;
    mem[121] = 8'h00;
    mem[122] = 8'h00;
    mem[123] = 8'h00;
    mem[124] = 8'h00;
    mem[125] = 8'h00;
    mem[126] = 8'h00;
    mem[127] = 8'h00;
    mem[128] = 8'h00;
    mem[129] = 8'h00;
    mem[130] = 8'h00;
    mem[131] = 8'h00;
    mem[132] = 8'h00;
    mem[133] = 8'h00;
    mem[134] = 8'h00;
    mem[135] = 8'h00;
    mem[136] = 8'h00;
    mem[137] = 8'h00;
    mem[138] = 8'hfc;
    mem[139] = 8'h00;
    mem[140] = 8'h00;
    mem[141] = 8'hfc;
    mem[142] = 8'h0f;
    mem[143] = 8'h00;
    mem[144] = 8'h00;
    mem[145] = 8'h00;
    mem[146] = 8'hff;
    mem[147] = 8'h00;
    mem[148] = 8'h00;
    mem[149] = 8'hff;
    mem[150] = 8'h1f;
    mem[151] = 8'h00;
    mem[152] = 8'h00;
    mem[153] = 8'h80;
    mem[154] = 8'hff;
    mem[155] = 8'h00;
    mem[156] = 8'h80;
    mem[157] = 8'hff;
    mem[158] = 8'h7f;
    mem[159] = 8'h00;
    mem[160] = 8'h00;
    mem[161] = 8'he0;
    mem[162] = 8'hff;
    mem[163] = 8'h00;
    mem[164] = 8'hc0;
    mem[165] = 8'h07;
    mem[166] = 8'h7c;
    mem[167] = 8'h00;
    mem[168] = 8'h00;
    mem[169] = 8'hf8;
    mem[170] = 8'hff;
    mem[171] = 8'h00;
    mem[172] = 8'he0;
    mem[173] = 8'h03;
    mem[174] = 8'hf8;
    mem[175] = 8'h00;
    mem[176] = 8'h00;
    mem[177] = 8'hfc;
    mem[178] = 8'hf9;
    mem[179] = 8'h00;
    mem[180] = 8'he0;
    mem[181] = 8'h01;
    mem[182] = 8'hf0;
    mem[183] = 8'h00;
    mem[184] = 8'h00;
    mem[185] = 8'h7c;
    mem[186] = 8'hf8;
    mem[187] = 8'h00;
    mem[188] = 8'hf0;
    mem[189] = 8'h00;
    mem[190] = 8'hf0;
    mem[191] = 8'h01;
    mem[192] = 8'h00;
    mem[193] = 8'h3c;
    mem[194] = 8'hf8;
    mem[195] = 8'h00;
    mem[196] = 8'hf0;
    mem[197] = 8'h00;
    mem[198] = 8'he0;
    mem[199] = 8'h01;
    mem[200] = 8'h00;
    mem[201] = 8'h0c;
    mem[202] = 8'hf8;
    mem[203] = 8'h00;
    mem[204] = 8'h78;
    mem[205] = 8'h00;
    mem[206] = 8'he0;
    mem[207] = 8'h01;
    mem[208] = 8'h00;
    mem[209] = 8'h00;
    mem[210] = 8'hf8;
    mem[211] = 8'h00;
    mem[212] = 8'h78;
    mem[213] = 8'h00;
    mem[214] = 8'h00;
    mem[215] = 8'h00;
    mem[216] = 8'h00;
    mem[217] = 8'h00;
    mem[218] = 8'hf8;
    mem[219] = 8'h00;
    mem[220] = 8'h78;
    mem[221] = 8'h00;
    mem[222] = 8'h00;
    mem[223] = 8'h00;
    mem[224] = 8'h00;
    mem[225] = 8'h00;
    mem[226] = 8'hf8;
    mem[227] = 8'h00;
    mem[228] = 8'h78;
    mem[229] = 8'hf8;
    mem[230] = 8'h07;
    mem[231] = 8'h00;
    mem[232] = 8'h00;
    mem[233] = 8'h00;
    mem[234] = 8'hf8;
    mem[235] = 8'h00;
    mem[236] = 8'h7c;
    mem[237] = 8'hfe;
    mem[238] = 8'h1f;
    mem[239] = 8'h00;
    mem[240] = 8'h00;
    mem[241] = 8'h00;
    mem[242] = 8'hf8;
    mem[243] = 8'h00;
    mem[244] = 8'h7c;
    mem[245] = 8'hff;
    mem[246] = 8'h3f;
    mem[247] = 8'h00;
    mem[248] = 8'h00;
    mem[249] = 8'h00;
    mem[250] = 8'hf8;
    mem[251] = 8'h00;
    mem[252] = 8'hfc;
    mem[253] = 8'h07;
    mem[254] = 8'h7e;
    mem[255] = 8'h00;
    mem[256] = 8'h00;
    mem[257] = 8'h00;
    mem[258] = 8'hf8;
    mem[259] = 8'h00;
    mem[260] = 8'hfc;
    mem[261] = 8'h01;
    mem[262] = 8'hfc;
    mem[263] = 8'h00;
    mem[264] = 8'h00;
    mem[265] = 8'h00;
    mem[266] = 8'hf8;
    mem[267] = 8'h00;
    mem[268] = 8'hfc;
    mem[269] = 8'h00;
    mem[270] = 8'hf8;
    mem[271] = 8'h00;
    mem[272] = 8'h00;
    mem[273] = 8'h00;
    mem[274] = 8'hf8;
    mem[275] = 8'h00;
    mem[276] = 8'hfc;
    mem[277] = 8'h00;
    mem[278] = 8'hf0;
    mem[279] = 8'h01;
    mem[280] = 8'h00;
    mem[281] = 8'h00;
    mem[282] = 8'hf8;
    mem[283] = 8'h00;
    mem[284] = 8'h7c;
    mem[285] = 8'h00;
    mem[286] = 8'hf0;
    mem[287] = 8'h01;
    mem[288] = 8'h00;
    mem[289] = 8'h00;
    mem[290] = 8'hf8;
    mem[291] = 8'h00;
    mem[292] = 8'h7c;
    mem[293] = 8'h00;
    mem[294] = 8'he0;
    mem[295] = 8'h01;
    mem[296] = 8'h00;
    mem[297] = 8'h00;
    mem[298] = 8'hf8;
    mem[299] = 8'h00;
    mem[300] = 8'h7c;
    mem[301] = 8'h00;
    mem[302] = 8'he0;
    mem[303] = 8'h01;
    mem[304] = 8'h00;
    mem[305] = 8'h00;
    mem[306] = 8'hf8;
    mem[307] = 8'h00;
    mem[308] = 8'h7c;
    mem[309] = 8'h00;
    mem[310] = 8'he0;
    mem[311] = 8'h01;
    mem[312] = 8'h00;
    mem[313] = 8'h00;
    mem[314] = 8'hf8;
    mem[315] = 8'h00;
    mem[316] = 8'h7c;
    mem[317] = 8'h00;
    mem[318] = 8'he0;
    mem[319] = 8'h01;
    mem[320] = 8'h00;
    mem[321] = 8'h00;
    mem[322] = 8'hf8;
    mem[323] = 8'h00;
    mem[324] = 8'h7c;
    mem[325] = 8'h00;
    mem[326] = 8'he0;
    mem[327] = 8'h01;
    mem[328] = 8'h00;
    mem[329] = 8'h00;
    mem[330] = 8'hf8;
    mem[331] = 8'h00;
    mem[332] = 8'h78;
    mem[333] = 8'h00;
    mem[334] = 8'he0;
    mem[335] = 8'h01;
    mem[336] = 8'h00;
    mem[337] = 8'h00;
    mem[338] = 8'hf8;
    mem[339] = 8'h00;
    mem[340] = 8'h78;
    mem[341] = 8'h00;
    mem[342] = 8'hf0;
    mem[343] = 8'h01;
    mem[344] = 8'h00;
    mem[345] = 8'h00;
    mem[346] = 8'hf8;
    mem[347] = 8'h00;
    mem[348] = 8'h78;
    mem[349] = 8'h00;
    mem[350] = 8'hf0;
    mem[351] = 8'h01;
    mem[352] = 8'h00;
    mem[353] = 8'h00;
    mem[354] = 8'hf8;
    mem[355] = 8'h00;
    mem[356] = 8'hf0;
    mem[357] = 8'h00;
    mem[358] = 8'hf8;
    mem[359] = 8'h00;
    mem[360] = 8'h00;
    mem[361] = 8'h00;
    mem[362] = 8'hf8;
    mem[363] = 8'h00;
    mem[364] = 8'hf0;
    mem[365] = 8'h01;
    mem[366] = 8'hf8;
    mem[367] = 8'h00;
    mem[368] = 8'h00;
    mem[369] = 8'h00;
    mem[370] = 8'hf8;
    mem[371] = 8'h00;
    mem[372] = 8'he0;
    mem[373] = 8'h03;
    mem[374] = 8'h7e;
    mem[375] = 8'h00;
    mem[376] = 8'h00;
    mem[377] = 8'h00;
    mem[378] = 8'hf8;
    mem[379] = 8'h00;
    mem[380] = 8'hc0;
    mem[381] = 8'hff;
    mem[382] = 8'h3f;
    mem[383] = 8'h00;
    mem[384] = 8'h00;
    mem[385] = 8'h00;
    mem[386] = 8'hf8;
    mem[387] = 8'h00;
    mem[388] = 8'h80;
    mem[389] = 8'hff;
    mem[390] = 8'h1f;
    mem[391] = 8'h00;
    mem[392] = 8'h00;
    mem[393] = 8'h00;
    mem[394] = 8'hf8;
    mem[395] = 8'h00;
    mem[396] = 8'h00;
    mem[397] = 8'hfe;
    mem[398] = 8'h07;
    mem[399] = 8'h00;
    mem[400] = 8'h00;
    mem[401] = 8'h00;
    mem[402] = 8'h00;
    mem[403] = 8'h00;
    mem[404] = 8'h00;
    mem[405] = 8'h00;
    mem[406] = 8'h00;
    mem[407] = 8'h00;
    mem[408] = 8'h00;
    mem[409] = 8'h00;
    mem[410] = 8'h00;
    mem[411] = 8'h00;
    mem[412] = 8'h00;
    mem[413] = 8'h00;
    mem[414] = 8'h00;
    mem[415] = 8'h00;
    mem[416] = 8'h00;
    mem[417] = 8'h00;
    mem[418] = 8'h00;
    mem[419] = 8'h00;
    mem[420] = 8'h00;
    mem[421] = 8'h00;
    mem[422] = 8'h00;
    mem[423] = 8'h00;
    mem[424] = 8'h00;
    mem[425] = 8'h00;
    mem[426] = 8'h00;
    mem[427] = 8'h00;
    mem[428] = 8'h00;
    mem[429] = 8'h00;
    mem[430] = 8'h00;
    mem[431] = 8'h00;
    mem[432] = 8'h00;
    mem[433] = 8'h00;
    mem[434] = 8'h00;
    mem[435] = 8'h00;
    mem[436] = 8'h00;
    mem[437] = 8'h00;
    mem[438] = 8'h00;
    mem[439] = 8'h00;
    mem[440] = 8'h00;
    mem[441] = 8'h00;
    mem[442] = 8'h00;
    mem[443] = 8'h00;
    mem[444] = 8'h00;
    mem[445] = 8'h00;
    mem[446] = 8'h00;
    mem[447] = 8'h00;
    mem[448] = 8'h00;
    mem[449] = 8'h00;
    mem[450] = 8'h00;
    mem[451] = 8'h00;
    mem[452] = 8'h00;
    mem[453] = 8'h00;
    mem[454] = 8'h00;
    mem[455] = 8'h00;
    mem[456] = 8'h00;
    mem[457] = 8'h00;
    mem[458] = 8'h00;
    mem[459] = 8'h00;
    mem[460] = 8'h00;
    mem[461] = 8'h00;
    mem[462] = 8'h00;
    mem[463] = 8'h00;
    mem[464] = 8'h00;
    mem[465] = 8'h00;
    mem[466] = 8'h00;
    mem[467] = 8'h00;
    mem[468] = 8'h00;
    mem[469] = 8'h00;
    mem[470] = 8'h00;
    mem[471] = 8'h00;
    mem[472] = 8'h00;
    mem[473] = 8'h00;
    mem[474] = 8'h00;
    mem[475] = 8'h00;
    mem[476] = 8'h00;
    mem[477] = 8'h00;
    mem[478] = 8'h00;
    mem[479] = 8'h00;
    mem[480] = 8'h00;
    mem[481] = 8'h00;
    mem[482] = 8'h00;
    mem[483] = 8'h00;
    mem[484] = 8'h00;
    mem[485] = 8'h00;
    mem[486] = 8'h00;
    mem[487] = 8'h00;
    mem[488] = 8'h00;
    mem[489] = 8'h00;
    mem[490] = 8'h00;
    mem[491] = 8'h00;
    mem[492] = 8'h00;
    mem[493] = 8'h00;
    mem[494] = 8'h00;
    mem[495] = 8'h00;
    mem[496] = 8'h00;
    mem[497] = 8'h00;
    mem[498] = 8'h00;
    mem[499] = 8'h00;
    mem[500] = 8'h00;
    mem[501] = 8'h00;
    mem[502] = 8'h00;
    mem[503] = 8'h00;
    mem[504] = 8'h00;
    mem[505] = 8'h00;
    mem[506] = 8'h00;
    mem[507] = 8'h00;
    mem[508] = 8'h00;
    mem[509] = 8'h00;
    mem[510] = 8'h00;
    mem[511] = 8'h00;
  end

  wire [8:0] addr = {y[5:0], x[5:3]};
  assign pixel = mem[addr][x&7];

endmodule

module glyph_32 (
    input wire [5:0] x,
    input wire [5:0] y,
    output wire pixel
);

  reg [7:0] mem[511:0];
  initial begin
    mem[0] = 8'h00;
    mem[1] = 8'h00;
    mem[2] = 8'h00;
    mem[3] = 8'h00;
    mem[4] = 8'h00;
    mem[5] = 8'h00;
    mem[6] = 8'h00;
    mem[7] = 8'h00;
    mem[8] = 8'h00;
    mem[9] = 8'h00;
    mem[10] = 8'h00;
    mem[11] = 8'h00;
    mem[12] = 8'h00;
    mem[13] = 8'h00;
    mem[14] = 8'h00;
    mem[15] = 8'h00;
    mem[16] = 8'h00;
    mem[17] = 8'h00;
    mem[18] = 8'h00;
    mem[19] = 8'h00;
    mem[20] = 8'h00;
    mem[21] = 8'h00;
    mem[22] = 8'h00;
    mem[23] = 8'h00;
    mem[24] = 8'h00;
    mem[25] = 8'h00;
    mem[26] = 8'h00;
    mem[27] = 8'h00;
    mem[28] = 8'h00;
    mem[29] = 8'h00;
    mem[30] = 8'h00;
    mem[31] = 8'h00;
    mem[32] = 8'h00;
    mem[33] = 8'h00;
    mem[34] = 8'h00;
    mem[35] = 8'h00;
    mem[36] = 8'h00;
    mem[37] = 8'h00;
    mem[38] = 8'h00;
    mem[39] = 8'h00;
    mem[40] = 8'h00;
    mem[41] = 8'h00;
    mem[42] = 8'h00;
    mem[43] = 8'h00;
    mem[44] = 8'h00;
    mem[45] = 8'h00;
    mem[46] = 8'h00;
    mem[47] = 8'h00;
    mem[48] = 8'h00;
    mem[49] = 8'h00;
    mem[50] = 8'h00;
    mem[51] = 8'h00;
    mem[52] = 8'h00;
    mem[53] = 8'h00;
    mem[54] = 8'h00;
    mem[55] = 8'h00;
    mem[56] = 8'h00;
    mem[57] = 8'h00;
    mem[58] = 8'h00;
    mem[59] = 8'h00;
    mem[60] = 8'h00;
    mem[61] = 8'h00;
    mem[62] = 8'h00;
    mem[63] = 8'h00;
    mem[64] = 8'h00;
    mem[65] = 8'h00;
    mem[66] = 8'h00;
    mem[67] = 8'h00;
    mem[68] = 8'h00;
    mem[69] = 8'h00;
    mem[70] = 8'h00;
    mem[71] = 8'h00;
    mem[72] = 8'h00;
    mem[73] = 8'h00;
    mem[74] = 8'h00;
    mem[75] = 8'h00;
    mem[76] = 8'h00;
    mem[77] = 8'h00;
    mem[78] = 8'h00;
    mem[79] = 8'h00;
    mem[80] = 8'h00;
    mem[81] = 8'h00;
    mem[82] = 8'h00;
    mem[83] = 8'h00;
    mem[84] = 8'h00;
    mem[85] = 8'h00;
    mem[86] = 8'h00;
    mem[87] = 8'h00;
    mem[88] = 8'h00;
    mem[89] = 8'h00;
    mem[90] = 8'h00;
    mem[91] = 8'h00;
    mem[92] = 8'h00;
    mem[93] = 8'h00;
    mem[94] = 8'h00;
    mem[95] = 8'h00;
    mem[96] = 8'h00;
    mem[97] = 8'h00;
    mem[98] = 8'h00;
    mem[99] = 8'h00;
    mem[100] = 8'h00;
    mem[101] = 8'h00;
    mem[102] = 8'h00;
    mem[103] = 8'h00;
    mem[104] = 8'h00;
    mem[105] = 8'h00;
    mem[106] = 8'h00;
    mem[107] = 8'h00;
    mem[108] = 8'h00;
    mem[109] = 8'h00;
    mem[110] = 8'h00;
    mem[111] = 8'h00;
    mem[112] = 8'h00;
    mem[113] = 8'h00;
    mem[114] = 8'h00;
    mem[115] = 8'h00;
    mem[116] = 8'h00;
    mem[117] = 8'h00;
    mem[118] = 8'h00;
    mem[119] = 8'h00;
    mem[120] = 8'h00;
    mem[121] = 8'h00;
    mem[122] = 8'h00;
    mem[123] = 8'h00;
    mem[124] = 8'h00;
    mem[125] = 8'h00;
    mem[126] = 8'h00;
    mem[127] = 8'h00;
    mem[128] = 8'h00;
    mem[129] = 8'h00;
    mem[130] = 8'h00;
    mem[131] = 8'h00;
    mem[132] = 8'h00;
    mem[133] = 8'h00;
    mem[134] = 8'h00;
    mem[135] = 8'h00;
    mem[136] = 8'h00;
    mem[137] = 8'he0;
    mem[138] = 8'hff;
    mem[139] = 8'h00;
    mem[140] = 8'h00;
    mem[141] = 8'hfc;
    mem[142] = 8'h0f;
    mem[143] = 8'h00;
    mem[144] = 8'h00;
    mem[145] = 8'hf8;
    mem[146] = 8'hff;
    mem[147] = 8'h01;
    mem[148] = 8'h00;
    mem[149] = 8'hff;
    mem[150] = 8'h3f;
    mem[151] = 8'h00;
    mem[152] = 8'h00;
    mem[153] = 8'hfc;
    mem[154] = 8'hff;
    mem[155] = 8'h07;
    mem[156] = 8'h80;
    mem[157] = 8'hff;
    mem[158] = 8'h7f;
    mem[159] = 8'h00;
    mem[160] = 8'h00;
    mem[161] = 8'h7e;
    mem[162] = 8'he0;
    mem[163] = 8'h07;
    mem[164] = 8'hc0;
    mem[165] = 8'h07;
    mem[166] = 8'hfc;
    mem[167] = 8'h00;
    mem[168] = 8'h00;
    mem[169] = 8'h1e;
    mem[170] = 8'h80;
    mem[171] = 8'h0f;
    mem[172] = 8'hc0;
    mem[173] = 8'h03;
    mem[174] = 8'hf8;
    mem[175] = 8'h01;
    mem[176] = 8'h00;
    mem[177] = 8'h1f;
    mem[178] = 8'h80;
    mem[179] = 8'h0f;
    mem[180] = 8'he0;
    mem[181] = 8'h01;
    mem[182] = 8'hf0;
    mem[183] = 8'h01;
    mem[184] = 8'h00;
    mem[185] = 8'h0f;
    mem[186] = 8'h00;
    mem[187] = 8'h0f;
    mem[188] = 8'he0;
    mem[189] = 8'h01;
    mem[190] = 8'he0;
    mem[191] = 8'h01;
    mem[192] = 8'h80;
    mem[193] = 8'h0f;
    mem[194] = 8'h00;
    mem[195] = 8'h0f;
    mem[196] = 8'hf0;
    mem[197] = 8'h01;
    mem[198] = 8'he0;
    mem[199] = 8'h01;
    mem[200] = 8'h80;
    mem[201] = 8'h07;
    mem[202] = 8'h00;
    mem[203] = 8'h0f;
    mem[204] = 8'hf0;
    mem[205] = 8'h00;
    mem[206] = 8'he0;
    mem[207] = 8'h01;
    mem[208] = 8'h80;
    mem[209] = 8'h07;
    mem[210] = 8'h00;
    mem[211] = 8'h0f;
    mem[212] = 8'hf0;
    mem[213] = 8'h00;
    mem[214] = 8'he0;
    mem[215] = 8'h01;
    mem[216] = 8'h00;
    mem[217] = 8'h00;
    mem[218] = 8'h00;
    mem[219] = 8'h0f;
    mem[220] = 8'h00;
    mem[221] = 8'h00;
    mem[222] = 8'he0;
    mem[223] = 8'h01;
    mem[224] = 8'h00;
    mem[225] = 8'h00;
    mem[226] = 8'h80;
    mem[227] = 8'h0f;
    mem[228] = 8'h00;
    mem[229] = 8'h00;
    mem[230] = 8'he0;
    mem[231] = 8'h01;
    mem[232] = 8'h00;
    mem[233] = 8'h00;
    mem[234] = 8'h80;
    mem[235] = 8'h07;
    mem[236] = 8'h00;
    mem[237] = 8'h00;
    mem[238] = 8'hf0;
    mem[239] = 8'h01;
    mem[240] = 8'h00;
    mem[241] = 8'h00;
    mem[242] = 8'he0;
    mem[243] = 8'h03;
    mem[244] = 8'h00;
    mem[245] = 8'h00;
    mem[246] = 8'hf0;
    mem[247] = 8'h00;
    mem[248] = 8'h00;
    mem[249] = 8'h00;
    mem[250] = 8'hf8;
    mem[251] = 8'h01;
    mem[252] = 8'h00;
    mem[253] = 8'h00;
    mem[254] = 8'hf8;
    mem[255] = 8'h00;
    mem[256] = 8'h00;
    mem[257] = 8'h00;
    mem[258] = 8'h7f;
    mem[259] = 8'h00;
    mem[260] = 8'h00;
    mem[261] = 8'h00;
    mem[262] = 8'h7c;
    mem[263] = 8'h00;
    mem[264] = 8'h00;
    mem[265] = 8'h00;
    mem[266] = 8'hff;
    mem[267] = 8'h01;
    mem[268] = 8'h00;
    mem[269] = 8'h00;
    mem[270] = 8'h3e;
    mem[271] = 8'h00;
    mem[272] = 8'h00;
    mem[273] = 8'h00;
    mem[274] = 8'hff;
    mem[275] = 8'h07;
    mem[276] = 8'h00;
    mem[277] = 8'h00;
    mem[278] = 8'h1f;
    mem[279] = 8'h00;
    mem[280] = 8'h00;
    mem[281] = 8'h00;
    mem[282] = 8'he0;
    mem[283] = 8'h0f;
    mem[284] = 8'h00;
    mem[285] = 8'h80;
    mem[286] = 8'h0f;
    mem[287] = 8'h00;
    mem[288] = 8'h00;
    mem[289] = 8'h00;
    mem[290] = 8'h80;
    mem[291] = 8'h0f;
    mem[292] = 8'h00;
    mem[293] = 8'hc0;
    mem[294] = 8'h0f;
    mem[295] = 8'h00;
    mem[296] = 8'h00;
    mem[297] = 8'h00;
    mem[298] = 8'h00;
    mem[299] = 8'h1f;
    mem[300] = 8'h00;
    mem[301] = 8'he0;
    mem[302] = 8'h07;
    mem[303] = 8'h00;
    mem[304] = 8'h00;
    mem[305] = 8'h00;
    mem[306] = 8'h00;
    mem[307] = 8'h1f;
    mem[308] = 8'h00;
    mem[309] = 8'hf0;
    mem[310] = 8'h03;
    mem[311] = 8'h00;
    mem[312] = 8'h00;
    mem[313] = 8'h00;
    mem[314] = 8'h00;
    mem[315] = 8'h1e;
    mem[316] = 8'h00;
    mem[317] = 8'hf8;
    mem[318] = 8'h01;
    mem[319] = 8'h00;
    mem[320] = 8'hc0;
    mem[321] = 8'h03;
    mem[322] = 8'h00;
    mem[323] = 8'h1e;
    mem[324] = 8'h00;
    mem[325] = 8'hfc;
    mem[326] = 8'h00;
    mem[327] = 8'h00;
    mem[328] = 8'hc0;
    mem[329] = 8'h03;
    mem[330] = 8'h00;
    mem[331] = 8'h1e;
    mem[332] = 8'h00;
    mem[333] = 8'h7e;
    mem[334] = 8'h00;
    mem[335] = 8'h00;
    mem[336] = 8'hc0;
    mem[337] = 8'h03;
    mem[338] = 8'h00;
    mem[339] = 8'h1e;
    mem[340] = 8'h00;
    mem[341] = 8'h3f;
    mem[342] = 8'h00;
    mem[343] = 8'h00;
    mem[344] = 8'hc0;
    mem[345] = 8'h07;
    mem[346] = 8'h00;
    mem[347] = 8'h1e;
    mem[348] = 8'h80;
    mem[349] = 8'h0f;
    mem[350] = 8'h00;
    mem[351] = 8'h00;
    mem[352] = 8'h80;
    mem[353] = 8'h07;
    mem[354] = 8'h00;
    mem[355] = 8'h1f;
    mem[356] = 8'hc0;
    mem[357] = 8'h07;
    mem[358] = 8'h00;
    mem[359] = 8'h00;
    mem[360] = 8'h80;
    mem[361] = 8'h0f;
    mem[362] = 8'h80;
    mem[363] = 8'h0f;
    mem[364] = 8'he0;
    mem[365] = 8'h03;
    mem[366] = 8'h00;
    mem[367] = 8'h00;
    mem[368] = 8'h00;
    mem[369] = 8'h3f;
    mem[370] = 8'hc0;
    mem[371] = 8'h07;
    mem[372] = 8'hf0;
    mem[373] = 8'h03;
    mem[374] = 8'h00;
    mem[375] = 8'h00;
    mem[376] = 8'h00;
    mem[377] = 8'hfe;
    mem[378] = 8'hff;
    mem[379] = 8'h03;
    mem[380] = 8'hf8;
    mem[381] = 8'hff;
    mem[382] = 8'hff;
    mem[383] = 8'h03;
    mem[384] = 8'h00;
    mem[385] = 8'hfc;
    mem[386] = 8'hff;
    mem[387] = 8'h01;
    mem[388] = 8'hf8;
    mem[389] = 8'hff;
    mem[390] = 8'hff;
    mem[391] = 8'h03;
    mem[392] = 8'h00;
    mem[393] = 8'hf0;
    mem[394] = 8'h7f;
    mem[395] = 8'h00;
    mem[396] = 8'hf8;
    mem[397] = 8'hff;
    mem[398] = 8'hff;
    mem[399] = 8'h03;
    mem[400] = 8'h00;
    mem[401] = 8'h00;
    mem[402] = 8'h00;
    mem[403] = 8'h00;
    mem[404] = 8'h00;
    mem[405] = 8'h00;
    mem[406] = 8'h00;
    mem[407] = 8'h00;
    mem[408] = 8'h00;
    mem[409] = 8'h00;
    mem[410] = 8'h00;
    mem[411] = 8'h00;
    mem[412] = 8'h00;
    mem[413] = 8'h00;
    mem[414] = 8'h00;
    mem[415] = 8'h00;
    mem[416] = 8'h00;
    mem[417] = 8'h00;
    mem[418] = 8'h00;
    mem[419] = 8'h00;
    mem[420] = 8'h00;
    mem[421] = 8'h00;
    mem[422] = 8'h00;
    mem[423] = 8'h00;
    mem[424] = 8'h00;
    mem[425] = 8'h00;
    mem[426] = 8'h00;
    mem[427] = 8'h00;
    mem[428] = 8'h00;
    mem[429] = 8'h00;
    mem[430] = 8'h00;
    mem[431] = 8'h00;
    mem[432] = 8'h00;
    mem[433] = 8'h00;
    mem[434] = 8'h00;
    mem[435] = 8'h00;
    mem[436] = 8'h00;
    mem[437] = 8'h00;
    mem[438] = 8'h00;
    mem[439] = 8'h00;
    mem[440] = 8'h00;
    mem[441] = 8'h00;
    mem[442] = 8'h00;
    mem[443] = 8'h00;
    mem[444] = 8'h00;
    mem[445] = 8'h00;
    mem[446] = 8'h00;
    mem[447] = 8'h00;
    mem[448] = 8'h00;
    mem[449] = 8'h00;
    mem[450] = 8'h00;
    mem[451] = 8'h00;
    mem[452] = 8'h00;
    mem[453] = 8'h00;
    mem[454] = 8'h00;
    mem[455] = 8'h00;
    mem[456] = 8'h00;
    mem[457] = 8'h00;
    mem[458] = 8'h00;
    mem[459] = 8'h00;
    mem[460] = 8'h00;
    mem[461] = 8'h00;
    mem[462] = 8'h00;
    mem[463] = 8'h00;
    mem[464] = 8'h00;
    mem[465] = 8'h00;
    mem[466] = 8'h00;
    mem[467] = 8'h00;
    mem[468] = 8'h00;
    mem[469] = 8'h00;
    mem[470] = 8'h00;
    mem[471] = 8'h00;
    mem[472] = 8'h00;
    mem[473] = 8'h00;
    mem[474] = 8'h00;
    mem[475] = 8'h00;
    mem[476] = 8'h00;
    mem[477] = 8'h00;
    mem[478] = 8'h00;
    mem[479] = 8'h00;
    mem[480] = 8'h00;
    mem[481] = 8'h00;
    mem[482] = 8'h00;
    mem[483] = 8'h00;
    mem[484] = 8'h00;
    mem[485] = 8'h00;
    mem[486] = 8'h00;
    mem[487] = 8'h00;
    mem[488] = 8'h00;
    mem[489] = 8'h00;
    mem[490] = 8'h00;
    mem[491] = 8'h00;
    mem[492] = 8'h00;
    mem[493] = 8'h00;
    mem[494] = 8'h00;
    mem[495] = 8'h00;
    mem[496] = 8'h00;
    mem[497] = 8'h00;
    mem[498] = 8'h00;
    mem[499] = 8'h00;
    mem[500] = 8'h00;
    mem[501] = 8'h00;
    mem[502] = 8'h00;
    mem[503] = 8'h00;
    mem[504] = 8'h00;
    mem[505] = 8'h00;
    mem[506] = 8'h00;
    mem[507] = 8'h00;
    mem[508] = 8'h00;
    mem[509] = 8'h00;
    mem[510] = 8'h00;
    mem[511] = 8'h00;
  end

  wire [8:0] addr = {y[5:0], x[5:3]};
  assign pixel = mem[addr][x&7];

endmodule

module glyph_64 (
    input wire [5:0] x,
    input wire [5:0] y,
    output wire pixel
);

  reg [7:0] mem[511:0];
  initial begin
    mem[0] = 8'h00;
    mem[1] = 8'h00;
    mem[2] = 8'h00;
    mem[3] = 8'h00;
    mem[4] = 8'h00;
    mem[5] = 8'h00;
    mem[6] = 8'h00;
    mem[7] = 8'h00;
    mem[8] = 8'h00;
    mem[9] = 8'h00;
    mem[10] = 8'h00;
    mem[11] = 8'h00;
    mem[12] = 8'h00;
    mem[13] = 8'h00;
    mem[14] = 8'h00;
    mem[15] = 8'h00;
    mem[16] = 8'h00;
    mem[17] = 8'h00;
    mem[18] = 8'h00;
    mem[19] = 8'h00;
    mem[20] = 8'h00;
    mem[21] = 8'h00;
    mem[22] = 8'h00;
    mem[23] = 8'h00;
    mem[24] = 8'h00;
    mem[25] = 8'h00;
    mem[26] = 8'h00;
    mem[27] = 8'h00;
    mem[28] = 8'h00;
    mem[29] = 8'h00;
    mem[30] = 8'h00;
    mem[31] = 8'h00;
    mem[32] = 8'h00;
    mem[33] = 8'h00;
    mem[34] = 8'h00;
    mem[35] = 8'h00;
    mem[36] = 8'h00;
    mem[37] = 8'h00;
    mem[38] = 8'h00;
    mem[39] = 8'h00;
    mem[40] = 8'h00;
    mem[41] = 8'h00;
    mem[42] = 8'h00;
    mem[43] = 8'h00;
    mem[44] = 8'h00;
    mem[45] = 8'h00;
    mem[46] = 8'h00;
    mem[47] = 8'h00;
    mem[48] = 8'h00;
    mem[49] = 8'h00;
    mem[50] = 8'h00;
    mem[51] = 8'h00;
    mem[52] = 8'h00;
    mem[53] = 8'h00;
    mem[54] = 8'h00;
    mem[55] = 8'h00;
    mem[56] = 8'h00;
    mem[57] = 8'h00;
    mem[58] = 8'h00;
    mem[59] = 8'h00;
    mem[60] = 8'h00;
    mem[61] = 8'h00;
    mem[62] = 8'h00;
    mem[63] = 8'h00;
    mem[64] = 8'h00;
    mem[65] = 8'h00;
    mem[66] = 8'h00;
    mem[67] = 8'h00;
    mem[68] = 8'h00;
    mem[69] = 8'h00;
    mem[70] = 8'h00;
    mem[71] = 8'h00;
    mem[72] = 8'h00;
    mem[73] = 8'h00;
    mem[74] = 8'h00;
    mem[75] = 8'h00;
    mem[76] = 8'h00;
    mem[77] = 8'h00;
    mem[78] = 8'h00;
    mem[79] = 8'h00;
    mem[80] = 8'h00;
    mem[81] = 8'h00;
    mem[82] = 8'h00;
    mem[83] = 8'h00;
    mem[84] = 8'h00;
    mem[85] = 8'h00;
    mem[86] = 8'h00;
    mem[87] = 8'h00;
    mem[88] = 8'h00;
    mem[89] = 8'h00;
    mem[90] = 8'h00;
    mem[91] = 8'h00;
    mem[92] = 8'h00;
    mem[93] = 8'h00;
    mem[94] = 8'h00;
    mem[95] = 8'h00;
    mem[96] = 8'h00;
    mem[97] = 8'h00;
    mem[98] = 8'h00;
    mem[99] = 8'h00;
    mem[100] = 8'h00;
    mem[101] = 8'h00;
    mem[102] = 8'h00;
    mem[103] = 8'h00;
    mem[104] = 8'h00;
    mem[105] = 8'h00;
    mem[106] = 8'h00;
    mem[107] = 8'h00;
    mem[108] = 8'h00;
    mem[109] = 8'h00;
    mem[110] = 8'h00;
    mem[111] = 8'h00;
    mem[112] = 8'h00;
    mem[113] = 8'h00;
    mem[114] = 8'h00;
    mem[115] = 8'h00;
    mem[116] = 8'h00;
    mem[117] = 8'h00;
    mem[118] = 8'h00;
    mem[119] = 8'h00;
    mem[120] = 8'h00;
    mem[121] = 8'h00;
    mem[122] = 8'h00;
    mem[123] = 8'h00;
    mem[124] = 8'h00;
    mem[125] = 8'h00;
    mem[126] = 8'h00;
    mem[127] = 8'h00;
    mem[128] = 8'h00;
    mem[129] = 8'h00;
    mem[130] = 8'h00;
    mem[131] = 8'h00;
    mem[132] = 8'h00;
    mem[133] = 8'h00;
    mem[134] = 8'h00;
    mem[135] = 8'h00;
    mem[136] = 8'h00;
    mem[137] = 8'hc0;
    mem[138] = 8'hff;
    mem[139] = 8'h00;
    mem[140] = 8'h00;
    mem[141] = 8'h00;
    mem[142] = 8'h7c;
    mem[143] = 8'h00;
    mem[144] = 8'h00;
    mem[145] = 8'hf0;
    mem[146] = 8'hff;
    mem[147] = 8'h01;
    mem[148] = 8'h00;
    mem[149] = 8'h00;
    mem[150] = 8'h7e;
    mem[151] = 8'h00;
    mem[152] = 8'h00;
    mem[153] = 8'hf8;
    mem[154] = 8'hff;
    mem[155] = 8'h07;
    mem[156] = 8'h00;
    mem[157] = 8'h00;
    mem[158] = 8'h7f;
    mem[159] = 8'h00;
    mem[160] = 8'h00;
    mem[161] = 8'h7c;
    mem[162] = 8'hc0;
    mem[163] = 8'h07;
    mem[164] = 8'h00;
    mem[165] = 8'h00;
    mem[166] = 8'h7f;
    mem[167] = 8'h00;
    mem[168] = 8'h00;
    mem[169] = 8'h3e;
    mem[170] = 8'h80;
    mem[171] = 8'h0f;
    mem[172] = 8'h00;
    mem[173] = 8'h80;
    mem[174] = 8'h7f;
    mem[175] = 8'h00;
    mem[176] = 8'h00;
    mem[177] = 8'h1e;
    mem[178] = 8'h00;
    mem[179] = 8'h0f;
    mem[180] = 8'h00;
    mem[181] = 8'hc0;
    mem[182] = 8'h7f;
    mem[183] = 8'h00;
    mem[184] = 8'h00;
    mem[185] = 8'h0f;
    mem[186] = 8'h00;
    mem[187] = 8'h1f;
    mem[188] = 8'h00;
    mem[189] = 8'he0;
    mem[190] = 8'h7d;
    mem[191] = 8'h00;
    mem[192] = 8'h00;
    mem[193] = 8'h0f;
    mem[194] = 8'h00;
    mem[195] = 8'h1e;
    mem[196] = 8'h00;
    mem[197] = 8'he0;
    mem[198] = 8'h7d;
    mem[199] = 8'h00;
    mem[200] = 8'h80;
    mem[201] = 8'h07;
    mem[202] = 8'h00;
    mem[203] = 8'h1e;
    mem[204] = 8'h00;
    mem[205] = 8'hf0;
    mem[206] = 8'h7c;
    mem[207] = 8'h00;
    mem[208] = 8'h80;
    mem[209] = 8'h07;
    mem[210] = 8'h00;
    mem[211] = 8'h00;
    mem[212] = 8'h00;
    mem[213] = 8'hf8;
    mem[214] = 8'h7c;
    mem[215] = 8'h00;
    mem[216] = 8'h80;
    mem[217] = 8'h07;
    mem[218] = 8'h00;
    mem[219] = 8'h00;
    mem[220] = 8'h00;
    mem[221] = 8'h78;
    mem[222] = 8'h7c;
    mem[223] = 8'h00;
    mem[224] = 8'h80;
    mem[225] = 8'h87;
    mem[226] = 8'h7f;
    mem[227] = 8'h00;
    mem[228] = 8'h00;
    mem[229] = 8'h3c;
    mem[230] = 8'h7c;
    mem[231] = 8'h00;
    mem[232] = 8'hc0;
    mem[233] = 8'he7;
    mem[234] = 8'hff;
    mem[235] = 8'h01;
    mem[236] = 8'h00;
    mem[237] = 8'h3e;
    mem[238] = 8'h7c;
    mem[239] = 8'h00;
    mem[240] = 8'hc0;
    mem[241] = 8'hf7;
    mem[242] = 8'hff;
    mem[243] = 8'h03;
    mem[244] = 8'h00;
    mem[245] = 8'h1e;
    mem[246] = 8'h7c;
    mem[247] = 8'h00;
    mem[248] = 8'hc0;
    mem[249] = 8'h7f;
    mem[250] = 8'he0;
    mem[251] = 8'h07;
    mem[252] = 8'h00;
    mem[253] = 8'h0f;
    mem[254] = 8'h7c;
    mem[255] = 8'h00;
    mem[256] = 8'hc0;
    mem[257] = 8'h1f;
    mem[258] = 8'hc0;
    mem[259] = 8'h0f;
    mem[260] = 8'h80;
    mem[261] = 8'h07;
    mem[262] = 8'h7c;
    mem[263] = 8'h00;
    mem[264] = 8'hc0;
    mem[265] = 8'h0f;
    mem[266] = 8'h80;
    mem[267] = 8'h0f;
    mem[268] = 8'h80;
    mem[269] = 8'h07;
    mem[270] = 8'h7c;
    mem[271] = 8'h00;
    mem[272] = 8'hc0;
    mem[273] = 8'h0f;
    mem[274] = 8'h00;
    mem[275] = 8'h1f;
    mem[276] = 8'hc0;
    mem[277] = 8'h03;
    mem[278] = 8'h7c;
    mem[279] = 8'h00;
    mem[280] = 8'hc0;
    mem[281] = 8'h07;
    mem[282] = 8'h00;
    mem[283] = 8'h1f;
    mem[284] = 8'he0;
    mem[285] = 8'h01;
    mem[286] = 8'h7c;
    mem[287] = 8'h00;
    mem[288] = 8'hc0;
    mem[289] = 8'h07;
    mem[290] = 8'h00;
    mem[291] = 8'h1e;
    mem[292] = 8'hf0;
    mem[293] = 8'h01;
    mem[294] = 8'h7c;
    mem[295] = 8'h00;
    mem[296] = 8'hc0;
    mem[297] = 8'h07;
    mem[298] = 8'h00;
    mem[299] = 8'h1e;
    mem[300] = 8'hf0;
    mem[301] = 8'h00;
    mem[302] = 8'h7c;
    mem[303] = 8'h00;
    mem[304] = 8'hc0;
    mem[305] = 8'h07;
    mem[306] = 8'h00;
    mem[307] = 8'h1e;
    mem[308] = 8'h78;
    mem[309] = 8'h00;
    mem[310] = 8'h7c;
    mem[311] = 8'h00;
    mem[312] = 8'hc0;
    mem[313] = 8'h07;
    mem[314] = 8'h00;
    mem[315] = 8'h1e;
    mem[316] = 8'hfc;
    mem[317] = 8'hff;
    mem[318] = 8'hff;
    mem[319] = 8'h07;
    mem[320] = 8'hc0;
    mem[321] = 8'h07;
    mem[322] = 8'h00;
    mem[323] = 8'h1e;
    mem[324] = 8'hfc;
    mem[325] = 8'hff;
    mem[326] = 8'hff;
    mem[327] = 8'h07;
    mem[328] = 8'h80;
    mem[329] = 8'h07;
    mem[330] = 8'h00;
    mem[331] = 8'h1e;
    mem[332] = 8'hfc;
    mem[333] = 8'hff;
    mem[334] = 8'hff;
    mem[335] = 8'h07;
    mem[336] = 8'h80;
    mem[337] = 8'h07;
    mem[338] = 8'h00;
    mem[339] = 8'h1f;
    mem[340] = 8'h00;
    mem[341] = 8'h00;
    mem[342] = 8'h7c;
    mem[343] = 8'h00;
    mem[344] = 8'h80;
    mem[345] = 8'h07;
    mem[346] = 8'h00;
    mem[347] = 8'h1f;
    mem[348] = 8'h00;
    mem[349] = 8'h00;
    mem[350] = 8'h7c;
    mem[351] = 8'h00;
    mem[352] = 8'h00;
    mem[353] = 8'h0f;
    mem[354] = 8'h80;
    mem[355] = 8'h0f;
    mem[356] = 8'h00;
    mem[357] = 8'h00;
    mem[358] = 8'h7c;
    mem[359] = 8'h00;
    mem[360] = 8'h00;
    mem[361] = 8'h1f;
    mem[362] = 8'h80;
    mem[363] = 8'h0f;
    mem[364] = 8'h00;
    mem[365] = 8'h00;
    mem[366] = 8'h7c;
    mem[367] = 8'h00;
    mem[368] = 8'h00;
    mem[369] = 8'h3e;
    mem[370] = 8'he0;
    mem[371] = 8'h07;
    mem[372] = 8'h00;
    mem[373] = 8'h00;
    mem[374] = 8'h7c;
    mem[375] = 8'h00;
    mem[376] = 8'h00;
    mem[377] = 8'hfc;
    mem[378] = 8'hff;
    mem[379] = 8'h03;
    mem[380] = 8'h00;
    mem[381] = 8'h00;
    mem[382] = 8'h7c;
    mem[383] = 8'h00;
    mem[384] = 8'h00;
    mem[385] = 8'hf8;
    mem[386] = 8'hff;
    mem[387] = 8'h01;
    mem[388] = 8'h00;
    mem[389] = 8'h00;
    mem[390] = 8'h7c;
    mem[391] = 8'h00;
    mem[392] = 8'h00;
    mem[393] = 8'he0;
    mem[394] = 8'h7f;
    mem[395] = 8'h00;
    mem[396] = 8'h00;
    mem[397] = 8'h00;
    mem[398] = 8'h7c;
    mem[399] = 8'h00;
    mem[400] = 8'h00;
    mem[401] = 8'h00;
    mem[402] = 8'h00;
    mem[403] = 8'h00;
    mem[404] = 8'h00;
    mem[405] = 8'h00;
    mem[406] = 8'h00;
    mem[407] = 8'h00;
    mem[408] = 8'h00;
    mem[409] = 8'h00;
    mem[410] = 8'h00;
    mem[411] = 8'h00;
    mem[412] = 8'h00;
    mem[413] = 8'h00;
    mem[414] = 8'h00;
    mem[415] = 8'h00;
    mem[416] = 8'h00;
    mem[417] = 8'h00;
    mem[418] = 8'h00;
    mem[419] = 8'h00;
    mem[420] = 8'h00;
    mem[421] = 8'h00;
    mem[422] = 8'h00;
    mem[423] = 8'h00;
    mem[424] = 8'h00;
    mem[425] = 8'h00;
    mem[426] = 8'h00;
    mem[427] = 8'h00;
    mem[428] = 8'h00;
    mem[429] = 8'h00;
    mem[430] = 8'h00;
    mem[431] = 8'h00;
    mem[432] = 8'h00;
    mem[433] = 8'h00;
    mem[434] = 8'h00;
    mem[435] = 8'h00;
    mem[436] = 8'h00;
    mem[437] = 8'h00;
    mem[438] = 8'h00;
    mem[439] = 8'h00;
    mem[440] = 8'h00;
    mem[441] = 8'h00;
    mem[442] = 8'h00;
    mem[443] = 8'h00;
    mem[444] = 8'h00;
    mem[445] = 8'h00;
    mem[446] = 8'h00;
    mem[447] = 8'h00;
    mem[448] = 8'h00;
    mem[449] = 8'h00;
    mem[450] = 8'h00;
    mem[451] = 8'h00;
    mem[452] = 8'h00;
    mem[453] = 8'h00;
    mem[454] = 8'h00;
    mem[455] = 8'h00;
    mem[456] = 8'h00;
    mem[457] = 8'h00;
    mem[458] = 8'h00;
    mem[459] = 8'h00;
    mem[460] = 8'h00;
    mem[461] = 8'h00;
    mem[462] = 8'h00;
    mem[463] = 8'h00;
    mem[464] = 8'h00;
    mem[465] = 8'h00;
    mem[466] = 8'h00;
    mem[467] = 8'h00;
    mem[468] = 8'h00;
    mem[469] = 8'h00;
    mem[470] = 8'h00;
    mem[471] = 8'h00;
    mem[472] = 8'h00;
    mem[473] = 8'h00;
    mem[474] = 8'h00;
    mem[475] = 8'h00;
    mem[476] = 8'h00;
    mem[477] = 8'h00;
    mem[478] = 8'h00;
    mem[479] = 8'h00;
    mem[480] = 8'h00;
    mem[481] = 8'h00;
    mem[482] = 8'h00;
    mem[483] = 8'h00;
    mem[484] = 8'h00;
    mem[485] = 8'h00;
    mem[486] = 8'h00;
    mem[487] = 8'h00;
    mem[488] = 8'h00;
    mem[489] = 8'h00;
    mem[490] = 8'h00;
    mem[491] = 8'h00;
    mem[492] = 8'h00;
    mem[493] = 8'h00;
    mem[494] = 8'h00;
    mem[495] = 8'h00;
    mem[496] = 8'h00;
    mem[497] = 8'h00;
    mem[498] = 8'h00;
    mem[499] = 8'h00;
    mem[500] = 8'h00;
    mem[501] = 8'h00;
    mem[502] = 8'h00;
    mem[503] = 8'h00;
    mem[504] = 8'h00;
    mem[505] = 8'h00;
    mem[506] = 8'h00;
    mem[507] = 8'h00;
    mem[508] = 8'h00;
    mem[509] = 8'h00;
    mem[510] = 8'h00;
    mem[511] = 8'h00;
  end

  wire [8:0] addr = {y[5:0], x[5:3]};
  assign pixel = mem[addr][x&7];

endmodule

module glyph_128 (
    input wire [5:0] x,
    input wire [5:0] y,
    output wire pixel
);

  reg [7:0] mem[511:0];
  initial begin
    mem[0] = 8'h00;
    mem[1] = 8'h00;
    mem[2] = 8'h00;
    mem[3] = 8'h00;
    mem[4] = 8'h00;
    mem[5] = 8'h00;
    mem[6] = 8'h00;
    mem[7] = 8'h00;
    mem[8] = 8'h00;
    mem[9] = 8'h00;
    mem[10] = 8'h00;
    mem[11] = 8'h00;
    mem[12] = 8'h00;
    mem[13] = 8'h00;
    mem[14] = 8'h00;
    mem[15] = 8'h00;
    mem[16] = 8'h00;
    mem[17] = 8'h00;
    mem[18] = 8'h00;
    mem[19] = 8'h00;
    mem[20] = 8'h00;
    mem[21] = 8'h00;
    mem[22] = 8'h00;
    mem[23] = 8'h00;
    mem[24] = 8'h00;
    mem[25] = 8'h00;
    mem[26] = 8'h00;
    mem[27] = 8'h00;
    mem[28] = 8'h00;
    mem[29] = 8'h00;
    mem[30] = 8'h00;
    mem[31] = 8'h00;
    mem[32] = 8'h00;
    mem[33] = 8'h00;
    mem[34] = 8'h00;
    mem[35] = 8'h00;
    mem[36] = 8'h00;
    mem[37] = 8'h00;
    mem[38] = 8'h00;
    mem[39] = 8'h00;
    mem[40] = 8'h00;
    mem[41] = 8'h00;
    mem[42] = 8'h00;
    mem[43] = 8'h00;
    mem[44] = 8'h00;
    mem[45] = 8'h00;
    mem[46] = 8'h00;
    mem[47] = 8'h00;
    mem[48] = 8'h00;
    mem[49] = 8'h00;
    mem[50] = 8'h00;
    mem[51] = 8'h00;
    mem[52] = 8'h00;
    mem[53] = 8'h00;
    mem[54] = 8'h00;
    mem[55] = 8'h00;
    mem[56] = 8'h00;
    mem[57] = 8'h00;
    mem[58] = 8'h00;
    mem[59] = 8'h00;
    mem[60] = 8'h00;
    mem[61] = 8'h00;
    mem[62] = 8'h00;
    mem[63] = 8'h00;
    mem[64] = 8'h00;
    mem[65] = 8'h00;
    mem[66] = 8'h00;
    mem[67] = 8'h00;
    mem[68] = 8'h00;
    mem[69] = 8'h00;
    mem[70] = 8'h00;
    mem[71] = 8'h00;
    mem[72] = 8'h00;
    mem[73] = 8'h00;
    mem[74] = 8'h00;
    mem[75] = 8'h00;
    mem[76] = 8'h00;
    mem[77] = 8'h00;
    mem[78] = 8'h00;
    mem[79] = 8'h00;
    mem[80] = 8'h00;
    mem[81] = 8'h00;
    mem[82] = 8'h00;
    mem[83] = 8'h00;
    mem[84] = 8'h00;
    mem[85] = 8'h00;
    mem[86] = 8'h00;
    mem[87] = 8'h00;
    mem[88] = 8'h00;
    mem[89] = 8'h00;
    mem[90] = 8'h00;
    mem[91] = 8'h00;
    mem[92] = 8'h00;
    mem[93] = 8'h00;
    mem[94] = 8'h00;
    mem[95] = 8'h00;
    mem[96] = 8'h00;
    mem[97] = 8'h00;
    mem[98] = 8'h00;
    mem[99] = 8'h00;
    mem[100] = 8'h00;
    mem[101] = 8'h00;
    mem[102] = 8'h00;
    mem[103] = 8'h00;
    mem[104] = 8'h00;
    mem[105] = 8'h00;
    mem[106] = 8'h00;
    mem[107] = 8'h00;
    mem[108] = 8'h00;
    mem[109] = 8'h00;
    mem[110] = 8'h00;
    mem[111] = 8'h00;
    mem[112] = 8'h00;
    mem[113] = 8'h00;
    mem[114] = 8'h00;
    mem[115] = 8'h00;
    mem[116] = 8'h00;
    mem[117] = 8'h00;
    mem[118] = 8'h00;
    mem[119] = 8'h00;
    mem[120] = 8'h00;
    mem[121] = 8'h00;
    mem[122] = 8'h00;
    mem[123] = 8'h00;
    mem[124] = 8'h00;
    mem[125] = 8'h00;
    mem[126] = 8'h00;
    mem[127] = 8'h00;
    mem[128] = 8'h00;
    mem[129] = 8'h00;
    mem[130] = 8'h00;
    mem[131] = 8'h00;
    mem[132] = 8'h00;
    mem[133] = 8'h00;
    mem[134] = 8'h00;
    mem[135] = 8'h00;
    mem[136] = 8'h00;
    mem[137] = 8'h00;
    mem[138] = 8'h00;
    mem[139] = 8'h00;
    mem[140] = 8'h00;
    mem[141] = 8'h00;
    mem[142] = 8'h00;
    mem[143] = 8'h00;
    mem[144] = 8'h00;
    mem[145] = 8'h00;
    mem[146] = 8'h00;
    mem[147] = 8'h00;
    mem[148] = 8'h00;
    mem[149] = 8'h00;
    mem[150] = 8'h00;
    mem[151] = 8'h00;
    mem[152] = 8'h00;
    mem[153] = 8'h00;
    mem[154] = 8'h00;
    mem[155] = 8'h00;
    mem[156] = 8'h00;
    mem[157] = 8'h00;
    mem[158] = 8'h00;
    mem[159] = 8'h00;
    mem[160] = 8'h00;
    mem[161] = 8'h78;
    mem[162] = 8'h00;
    mem[163] = 8'hf0;
    mem[164] = 8'h1f;
    mem[165] = 8'h00;
    mem[166] = 8'hff;
    mem[167] = 8'h03;
    mem[168] = 8'h00;
    mem[169] = 8'h7e;
    mem[170] = 8'h00;
    mem[171] = 8'hfc;
    mem[172] = 8'h3f;
    mem[173] = 8'h80;
    mem[174] = 8'hff;
    mem[175] = 8'h07;
    mem[176] = 8'h00;
    mem[177] = 8'h7f;
    mem[178] = 8'h00;
    mem[179] = 8'h3e;
    mem[180] = 8'h7c;
    mem[181] = 8'hc0;
    mem[182] = 8'h83;
    mem[183] = 8'h0f;
    mem[184] = 8'hc0;
    mem[185] = 8'h7f;
    mem[186] = 8'h00;
    mem[187] = 8'h0e;
    mem[188] = 8'h70;
    mem[189] = 8'hc0;
    mem[190] = 8'h01;
    mem[191] = 8'h0e;
    mem[192] = 8'he0;
    mem[193] = 8'h73;
    mem[194] = 8'h00;
    mem[195] = 8'h0f;
    mem[196] = 8'hf0;
    mem[197] = 8'he0;
    mem[198] = 8'h01;
    mem[199] = 8'h1e;
    mem[200] = 8'he0;
    mem[201] = 8'h70;
    mem[202] = 8'h00;
    mem[203] = 8'h07;
    mem[204] = 8'hf0;
    mem[205] = 8'he0;
    mem[206] = 8'h00;
    mem[207] = 8'h1c;
    mem[208] = 8'h60;
    mem[209] = 8'h70;
    mem[210] = 8'h00;
    mem[211] = 8'h07;
    mem[212] = 8'he0;
    mem[213] = 8'he0;
    mem[214] = 8'h00;
    mem[215] = 8'h1c;
    mem[216] = 8'h00;
    mem[217] = 8'h70;
    mem[218] = 8'h00;
    mem[219] = 8'h07;
    mem[220] = 8'hf0;
    mem[221] = 8'he0;
    mem[222] = 8'h01;
    mem[223] = 8'h1e;
    mem[224] = 8'h00;
    mem[225] = 8'h70;
    mem[226] = 8'h00;
    mem[227] = 8'h00;
    mem[228] = 8'hf0;
    mem[229] = 8'hc0;
    mem[230] = 8'h01;
    mem[231] = 8'h1e;
    mem[232] = 8'h00;
    mem[233] = 8'h70;
    mem[234] = 8'h00;
    mem[235] = 8'h00;
    mem[236] = 8'h70;
    mem[237] = 8'hc0;
    mem[238] = 8'h03;
    mem[239] = 8'h0f;
    mem[240] = 8'h00;
    mem[241] = 8'h70;
    mem[242] = 8'h00;
    mem[243] = 8'h00;
    mem[244] = 8'h78;
    mem[245] = 8'h80;
    mem[246] = 8'hcf;
    mem[247] = 8'h07;
    mem[248] = 8'h00;
    mem[249] = 8'h70;
    mem[250] = 8'h00;
    mem[251] = 8'h00;
    mem[252] = 8'h3c;
    mem[253] = 8'h00;
    mem[254] = 8'hff;
    mem[255] = 8'h01;
    mem[256] = 8'h00;
    mem[257] = 8'h70;
    mem[258] = 8'h00;
    mem[259] = 8'h00;
    mem[260] = 8'h1c;
    mem[261] = 8'h80;
    mem[262] = 8'hff;
    mem[263] = 8'h03;
    mem[264] = 8'h00;
    mem[265] = 8'h70;
    mem[266] = 8'h00;
    mem[267] = 8'h00;
    mem[268] = 8'h1e;
    mem[269] = 8'hc0;
    mem[270] = 8'h83;
    mem[271] = 8'h0f;
    mem[272] = 8'h00;
    mem[273] = 8'h70;
    mem[274] = 8'h00;
    mem[275] = 8'h00;
    mem[276] = 8'h0f;
    mem[277] = 8'he0;
    mem[278] = 8'h01;
    mem[279] = 8'h0e;
    mem[280] = 8'h00;
    mem[281] = 8'h70;
    mem[282] = 8'h00;
    mem[283] = 8'h80;
    mem[284] = 8'h07;
    mem[285] = 8'hf0;
    mem[286] = 8'h00;
    mem[287] = 8'h1e;
    mem[288] = 8'h00;
    mem[289] = 8'h70;
    mem[290] = 8'h00;
    mem[291] = 8'hc0;
    mem[292] = 8'h03;
    mem[293] = 8'hf0;
    mem[294] = 8'h00;
    mem[295] = 8'h1c;
    mem[296] = 8'h00;
    mem[297] = 8'h70;
    mem[298] = 8'h00;
    mem[299] = 8'he0;
    mem[300] = 8'h01;
    mem[301] = 8'h70;
    mem[302] = 8'h00;
    mem[303] = 8'h1c;
    mem[304] = 8'h00;
    mem[305] = 8'h70;
    mem[306] = 8'h00;
    mem[307] = 8'hf0;
    mem[308] = 8'h00;
    mem[309] = 8'h70;
    mem[310] = 8'h00;
    mem[311] = 8'h1c;
    mem[312] = 8'h00;
    mem[313] = 8'h70;
    mem[314] = 8'h00;
    mem[315] = 8'h78;
    mem[316] = 8'h00;
    mem[317] = 8'hf0;
    mem[318] = 8'h00;
    mem[319] = 8'h1c;
    mem[320] = 8'h00;
    mem[321] = 8'h70;
    mem[322] = 8'h00;
    mem[323] = 8'h3c;
    mem[324] = 8'h00;
    mem[325] = 8'hf0;
    mem[326] = 8'h00;
    mem[327] = 8'h1e;
    mem[328] = 8'h00;
    mem[329] = 8'h70;
    mem[330] = 8'h00;
    mem[331] = 8'h1e;
    mem[332] = 8'h00;
    mem[333] = 8'he0;
    mem[334] = 8'h01;
    mem[335] = 8'h1e;
    mem[336] = 8'h00;
    mem[337] = 8'h70;
    mem[338] = 8'h00;
    mem[339] = 8'h0f;
    mem[340] = 8'h00;
    mem[341] = 8'he0;
    mem[342] = 8'h03;
    mem[343] = 8'h0f;
    mem[344] = 8'h00;
    mem[345] = 8'h70;
    mem[346] = 8'h80;
    mem[347] = 8'hff;
    mem[348] = 8'hff;
    mem[349] = 8'hc0;
    mem[350] = 8'hff;
    mem[351] = 8'h07;
    mem[352] = 8'h00;
    mem[353] = 8'h70;
    mem[354] = 8'h80;
    mem[355] = 8'hff;
    mem[356] = 8'hff;
    mem[357] = 8'h00;
    mem[358] = 8'hff;
    mem[359] = 8'h01;
    mem[360] = 8'h00;
    mem[361] = 8'h00;
    mem[362] = 8'h00;
    mem[363] = 8'h00;
    mem[364] = 8'h00;
    mem[365] = 8'h00;
    mem[366] = 8'h00;
    mem[367] = 8'h00;
    mem[368] = 8'h00;
    mem[369] = 8'h00;
    mem[370] = 8'h00;
    mem[371] = 8'h00;
    mem[372] = 8'h00;
    mem[373] = 8'h00;
    mem[374] = 8'h00;
    mem[375] = 8'h00;
    mem[376] = 8'h00;
    mem[377] = 8'h00;
    mem[378] = 8'h00;
    mem[379] = 8'h00;
    mem[380] = 8'h00;
    mem[381] = 8'h00;
    mem[382] = 8'h00;
    mem[383] = 8'h00;
    mem[384] = 8'h00;
    mem[385] = 8'h00;
    mem[386] = 8'h00;
    mem[387] = 8'h00;
    mem[388] = 8'h00;
    mem[389] = 8'h00;
    mem[390] = 8'h00;
    mem[391] = 8'h00;
    mem[392] = 8'h00;
    mem[393] = 8'h00;
    mem[394] = 8'h00;
    mem[395] = 8'h00;
    mem[396] = 8'h00;
    mem[397] = 8'h00;
    mem[398] = 8'h00;
    mem[399] = 8'h00;
    mem[400] = 8'h00;
    mem[401] = 8'h00;
    mem[402] = 8'h00;
    mem[403] = 8'h00;
    mem[404] = 8'h00;
    mem[405] = 8'h00;
    mem[406] = 8'h00;
    mem[407] = 8'h00;
    mem[408] = 8'h00;
    mem[409] = 8'h00;
    mem[410] = 8'h00;
    mem[411] = 8'h00;
    mem[412] = 8'h00;
    mem[413] = 8'h00;
    mem[414] = 8'h00;
    mem[415] = 8'h00;
    mem[416] = 8'h00;
    mem[417] = 8'h00;
    mem[418] = 8'h00;
    mem[419] = 8'h00;
    mem[420] = 8'h00;
    mem[421] = 8'h00;
    mem[422] = 8'h00;
    mem[423] = 8'h00;
    mem[424] = 8'h00;
    mem[425] = 8'h00;
    mem[426] = 8'h00;
    mem[427] = 8'h00;
    mem[428] = 8'h00;
    mem[429] = 8'h00;
    mem[430] = 8'h00;
    mem[431] = 8'h00;
    mem[432] = 8'h00;
    mem[433] = 8'h00;
    mem[434] = 8'h00;
    mem[435] = 8'h00;
    mem[436] = 8'h00;
    mem[437] = 8'h00;
    mem[438] = 8'h00;
    mem[439] = 8'h00;
    mem[440] = 8'h00;
    mem[441] = 8'h00;
    mem[442] = 8'h00;
    mem[443] = 8'h00;
    mem[444] = 8'h00;
    mem[445] = 8'h00;
    mem[446] = 8'h00;
    mem[447] = 8'h00;
    mem[448] = 8'h00;
    mem[449] = 8'h00;
    mem[450] = 8'h00;
    mem[451] = 8'h00;
    mem[452] = 8'h00;
    mem[453] = 8'h00;
    mem[454] = 8'h00;
    mem[455] = 8'h00;
    mem[456] = 8'h00;
    mem[457] = 8'h00;
    mem[458] = 8'h00;
    mem[459] = 8'h00;
    mem[460] = 8'h00;
    mem[461] = 8'h00;
    mem[462] = 8'h00;
    mem[463] = 8'h00;
    mem[464] = 8'h00;
    mem[465] = 8'h00;
    mem[466] = 8'h00;
    mem[467] = 8'h00;
    mem[468] = 8'h00;
    mem[469] = 8'h00;
    mem[470] = 8'h00;
    mem[471] = 8'h00;
    mem[472] = 8'h00;
    mem[473] = 8'h00;
    mem[474] = 8'h00;
    mem[475] = 8'h00;
    mem[476] = 8'h00;
    mem[477] = 8'h00;
    mem[478] = 8'h00;
    mem[479] = 8'h00;
    mem[480] = 8'h00;
    mem[481] = 8'h00;
    mem[482] = 8'h00;
    mem[483] = 8'h00;
    mem[484] = 8'h00;
    mem[485] = 8'h00;
    mem[486] = 8'h00;
    mem[487] = 8'h00;
    mem[488] = 8'h00;
    mem[489] = 8'h00;
    mem[490] = 8'h00;
    mem[491] = 8'h00;
    mem[492] = 8'h00;
    mem[493] = 8'h00;
    mem[494] = 8'h00;
    mem[495] = 8'h00;
    mem[496] = 8'h00;
    mem[497] = 8'h00;
    mem[498] = 8'h00;
    mem[499] = 8'h00;
    mem[500] = 8'h00;
    mem[501] = 8'h00;
    mem[502] = 8'h00;
    mem[503] = 8'h00;
    mem[504] = 8'h00;
    mem[505] = 8'h00;
    mem[506] = 8'h00;
    mem[507] = 8'h00;
    mem[508] = 8'h00;
    mem[509] = 8'h00;
    mem[510] = 8'h00;
    mem[511] = 8'h00;
  end

  wire [8:0] addr = {y[5:0], x[5:3]};
  assign pixel = mem[addr][x&7];

endmodule

module glyph_256 (
    input wire [5:0] x,
    input wire [5:0] y,
    output wire pixel
);

  reg [7:0] mem[511:0];
  initial begin
    mem[0] = 8'h00;
    mem[1] = 8'h00;
    mem[2] = 8'h00;
    mem[3] = 8'h00;
    mem[4] = 8'h00;
    mem[5] = 8'h00;
    mem[6] = 8'h00;
    mem[7] = 8'h00;
    mem[8] = 8'h00;
    mem[9] = 8'h00;
    mem[10] = 8'h00;
    mem[11] = 8'h00;
    mem[12] = 8'h00;
    mem[13] = 8'h00;
    mem[14] = 8'h00;
    mem[15] = 8'h00;
    mem[16] = 8'h00;
    mem[17] = 8'h00;
    mem[18] = 8'h00;
    mem[19] = 8'h00;
    mem[20] = 8'h00;
    mem[21] = 8'h00;
    mem[22] = 8'h00;
    mem[23] = 8'h00;
    mem[24] = 8'h00;
    mem[25] = 8'h00;
    mem[26] = 8'h00;
    mem[27] = 8'h00;
    mem[28] = 8'h00;
    mem[29] = 8'h00;
    mem[30] = 8'h00;
    mem[31] = 8'h00;
    mem[32] = 8'h00;
    mem[33] = 8'h00;
    mem[34] = 8'h00;
    mem[35] = 8'h00;
    mem[36] = 8'h00;
    mem[37] = 8'h00;
    mem[38] = 8'h00;
    mem[39] = 8'h00;
    mem[40] = 8'h00;
    mem[41] = 8'h00;
    mem[42] = 8'h00;
    mem[43] = 8'h00;
    mem[44] = 8'h00;
    mem[45] = 8'h00;
    mem[46] = 8'h00;
    mem[47] = 8'h00;
    mem[48] = 8'h00;
    mem[49] = 8'h00;
    mem[50] = 8'h00;
    mem[51] = 8'h00;
    mem[52] = 8'h00;
    mem[53] = 8'h00;
    mem[54] = 8'h00;
    mem[55] = 8'h00;
    mem[56] = 8'h00;
    mem[57] = 8'h00;
    mem[58] = 8'h00;
    mem[59] = 8'h00;
    mem[60] = 8'h00;
    mem[61] = 8'h00;
    mem[62] = 8'h00;
    mem[63] = 8'h00;
    mem[64] = 8'h00;
    mem[65] = 8'h00;
    mem[66] = 8'h00;
    mem[67] = 8'h00;
    mem[68] = 8'h00;
    mem[69] = 8'h00;
    mem[70] = 8'h00;
    mem[71] = 8'h00;
    mem[72] = 8'h00;
    mem[73] = 8'h00;
    mem[74] = 8'h00;
    mem[75] = 8'h00;
    mem[76] = 8'h00;
    mem[77] = 8'h00;
    mem[78] = 8'h00;
    mem[79] = 8'h00;
    mem[80] = 8'h00;
    mem[81] = 8'h00;
    mem[82] = 8'h00;
    mem[83] = 8'h00;
    mem[84] = 8'h00;
    mem[85] = 8'h00;
    mem[86] = 8'h00;
    mem[87] = 8'h00;
    mem[88] = 8'h00;
    mem[89] = 8'h00;
    mem[90] = 8'h00;
    mem[91] = 8'h00;
    mem[92] = 8'h00;
    mem[93] = 8'h00;
    mem[94] = 8'h00;
    mem[95] = 8'h00;
    mem[96] = 8'h00;
    mem[97] = 8'h00;
    mem[98] = 8'h00;
    mem[99] = 8'h00;
    mem[100] = 8'h00;
    mem[101] = 8'h00;
    mem[102] = 8'h00;
    mem[103] = 8'h00;
    mem[104] = 8'h00;
    mem[105] = 8'h00;
    mem[106] = 8'h00;
    mem[107] = 8'h00;
    mem[108] = 8'h00;
    mem[109] = 8'h00;
    mem[110] = 8'h00;
    mem[111] = 8'h00;
    mem[112] = 8'h00;
    mem[113] = 8'h00;
    mem[114] = 8'h00;
    mem[115] = 8'h00;
    mem[116] = 8'h00;
    mem[117] = 8'h00;
    mem[118] = 8'h00;
    mem[119] = 8'h00;
    mem[120] = 8'h00;
    mem[121] = 8'h00;
    mem[122] = 8'h00;
    mem[123] = 8'h00;
    mem[124] = 8'h00;
    mem[125] = 8'h00;
    mem[126] = 8'h00;
    mem[127] = 8'h00;
    mem[128] = 8'h00;
    mem[129] = 8'h00;
    mem[130] = 8'h00;
    mem[131] = 8'h00;
    mem[132] = 8'h00;
    mem[133] = 8'h00;
    mem[134] = 8'h00;
    mem[135] = 8'h00;
    mem[136] = 8'h00;
    mem[137] = 8'h00;
    mem[138] = 8'h00;
    mem[139] = 8'h00;
    mem[140] = 8'h00;
    mem[141] = 8'h00;
    mem[142] = 8'h00;
    mem[143] = 8'h00;
    mem[144] = 8'h00;
    mem[145] = 8'h00;
    mem[146] = 8'h00;
    mem[147] = 8'h00;
    mem[148] = 8'h00;
    mem[149] = 8'h00;
    mem[150] = 8'h00;
    mem[151] = 8'h00;
    mem[152] = 8'h00;
    mem[153] = 8'h00;
    mem[154] = 8'h00;
    mem[155] = 8'h00;
    mem[156] = 8'h00;
    mem[157] = 8'h00;
    mem[158] = 8'h00;
    mem[159] = 8'h00;
    mem[160] = 8'h80;
    mem[161] = 8'hff;
    mem[162] = 8'h00;
    mem[163] = 8'hfe;
    mem[164] = 8'h7f;
    mem[165] = 8'h00;
    mem[166] = 8'hfc;
    mem[167] = 8'h03;
    mem[168] = 8'he0;
    mem[169] = 8'hff;
    mem[170] = 8'h01;
    mem[171] = 8'hfe;
    mem[172] = 8'h7f;
    mem[173] = 8'h00;
    mem[174] = 8'hff;
    mem[175] = 8'h07;
    mem[176] = 8'hf0;
    mem[177] = 8'he1;
    mem[178] = 8'h03;
    mem[179] = 8'h0e;
    mem[180] = 8'h00;
    mem[181] = 8'h80;
    mem[182] = 8'h87;
    mem[183] = 8'h0f;
    mem[184] = 8'h70;
    mem[185] = 8'h80;
    mem[186] = 8'h03;
    mem[187] = 8'h0e;
    mem[188] = 8'h00;
    mem[189] = 8'hc0;
    mem[190] = 8'h03;
    mem[191] = 8'h0e;
    mem[192] = 8'h78;
    mem[193] = 8'h80;
    mem[194] = 8'h07;
    mem[195] = 8'h0e;
    mem[196] = 8'h00;
    mem[197] = 8'hc0;
    mem[198] = 8'h01;
    mem[199] = 8'h1e;
    mem[200] = 8'h38;
    mem[201] = 8'h80;
    mem[202] = 8'h07;
    mem[203] = 8'h06;
    mem[204] = 8'h00;
    mem[205] = 8'he0;
    mem[206] = 8'h00;
    mem[207] = 8'h1c;
    mem[208] = 8'h38;
    mem[209] = 8'h00;
    mem[210] = 8'h07;
    mem[211] = 8'h06;
    mem[212] = 8'h00;
    mem[213] = 8'he0;
    mem[214] = 8'h00;
    mem[215] = 8'h1c;
    mem[216] = 8'h38;
    mem[217] = 8'h80;
    mem[218] = 8'h07;
    mem[219] = 8'h07;
    mem[220] = 8'h00;
    mem[221] = 8'he0;
    mem[222] = 8'h00;
    mem[223] = 8'h00;
    mem[224] = 8'h00;
    mem[225] = 8'h80;
    mem[226] = 8'h07;
    mem[227] = 8'he7;
    mem[228] = 8'h07;
    mem[229] = 8'hf0;
    mem[230] = 8'hf8;
    mem[231] = 8'h00;
    mem[232] = 8'h00;
    mem[233] = 8'h80;
    mem[234] = 8'h03;
    mem[235] = 8'hf7;
    mem[236] = 8'h1f;
    mem[237] = 8'h70;
    mem[238] = 8'hfe;
    mem[239] = 8'h03;
    mem[240] = 8'h00;
    mem[241] = 8'hc0;
    mem[242] = 8'h03;
    mem[243] = 8'h7f;
    mem[244] = 8'h3e;
    mem[245] = 8'h70;
    mem[246] = 8'hef;
    mem[247] = 8'h07;
    mem[248] = 8'h00;
    mem[249] = 8'he0;
    mem[250] = 8'h01;
    mem[251] = 8'h1f;
    mem[252] = 8'h78;
    mem[253] = 8'hf0;
    mem[254] = 8'h03;
    mem[255] = 8'h0f;
    mem[256] = 8'h00;
    mem[257] = 8'he0;
    mem[258] = 8'h00;
    mem[259] = 8'h0f;
    mem[260] = 8'hf0;
    mem[261] = 8'hf0;
    mem[262] = 8'h01;
    mem[263] = 8'h1e;
    mem[264] = 8'h00;
    mem[265] = 8'hf0;
    mem[266] = 8'h00;
    mem[267] = 8'h07;
    mem[268] = 8'hf0;
    mem[269] = 8'hf0;
    mem[270] = 8'h00;
    mem[271] = 8'h1e;
    mem[272] = 8'h00;
    mem[273] = 8'h78;
    mem[274] = 8'h00;
    mem[275] = 8'h00;
    mem[276] = 8'he0;
    mem[277] = 8'hf0;
    mem[278] = 8'h00;
    mem[279] = 8'h1c;
    mem[280] = 8'h00;
    mem[281] = 8'h3c;
    mem[282] = 8'h00;
    mem[283] = 8'h00;
    mem[284] = 8'he0;
    mem[285] = 8'h70;
    mem[286] = 8'h00;
    mem[287] = 8'h1c;
    mem[288] = 8'h00;
    mem[289] = 8'h1e;
    mem[290] = 8'h00;
    mem[291] = 8'h00;
    mem[292] = 8'he0;
    mem[293] = 8'h70;
    mem[294] = 8'h00;
    mem[295] = 8'h1c;
    mem[296] = 8'h00;
    mem[297] = 8'h0f;
    mem[298] = 8'h00;
    mem[299] = 8'h00;
    mem[300] = 8'he0;
    mem[301] = 8'h70;
    mem[302] = 8'h00;
    mem[303] = 8'h1c;
    mem[304] = 8'h80;
    mem[305] = 8'h07;
    mem[306] = 8'h80;
    mem[307] = 8'h03;
    mem[308] = 8'he0;
    mem[309] = 8'hf0;
    mem[310] = 8'h00;
    mem[311] = 8'h1c;
    mem[312] = 8'hc0;
    mem[313] = 8'h03;
    mem[314] = 8'h80;
    mem[315] = 8'h07;
    mem[316] = 8'he0;
    mem[317] = 8'he0;
    mem[318] = 8'h00;
    mem[319] = 8'h1c;
    mem[320] = 8'he0;
    mem[321] = 8'h01;
    mem[322] = 8'h00;
    mem[323] = 8'h07;
    mem[324] = 8'hf0;
    mem[325] = 8'he0;
    mem[326] = 8'h00;
    mem[327] = 8'h1e;
    mem[328] = 8'hf0;
    mem[329] = 8'h00;
    mem[330] = 8'h00;
    mem[331] = 8'h0f;
    mem[332] = 8'h78;
    mem[333] = 8'hc0;
    mem[334] = 8'h01;
    mem[335] = 8'h0f;
    mem[336] = 8'h78;
    mem[337] = 8'h00;
    mem[338] = 8'h00;
    mem[339] = 8'h1e;
    mem[340] = 8'h3c;
    mem[341] = 8'hc0;
    mem[342] = 8'h83;
    mem[343] = 8'h07;
    mem[344] = 8'hfc;
    mem[345] = 8'hff;
    mem[346] = 8'h07;
    mem[347] = 8'hfc;
    mem[348] = 8'h1f;
    mem[349] = 8'h80;
    mem[350] = 8'hff;
    mem[351] = 8'h03;
    mem[352] = 8'hfc;
    mem[353] = 8'hff;
    mem[354] = 8'h07;
    mem[355] = 8'hf8;
    mem[356] = 8'h0f;
    mem[357] = 8'h00;
    mem[358] = 8'hff;
    mem[359] = 8'h01;
    mem[360] = 8'h00;
    mem[361] = 8'h00;
    mem[362] = 8'h00;
    mem[363] = 8'h00;
    mem[364] = 8'h00;
    mem[365] = 8'h00;
    mem[366] = 8'h00;
    mem[367] = 8'h00;
    mem[368] = 8'h00;
    mem[369] = 8'h00;
    mem[370] = 8'h00;
    mem[371] = 8'h00;
    mem[372] = 8'h00;
    mem[373] = 8'h00;
    mem[374] = 8'h00;
    mem[375] = 8'h00;
    mem[376] = 8'h00;
    mem[377] = 8'h00;
    mem[378] = 8'h00;
    mem[379] = 8'h00;
    mem[380] = 8'h00;
    mem[381] = 8'h00;
    mem[382] = 8'h00;
    mem[383] = 8'h00;
    mem[384] = 8'h00;
    mem[385] = 8'h00;
    mem[386] = 8'h00;
    mem[387] = 8'h00;
    mem[388] = 8'h00;
    mem[389] = 8'h00;
    mem[390] = 8'h00;
    mem[391] = 8'h00;
    mem[392] = 8'h00;
    mem[393] = 8'h00;
    mem[394] = 8'h00;
    mem[395] = 8'h00;
    mem[396] = 8'h00;
    mem[397] = 8'h00;
    mem[398] = 8'h00;
    mem[399] = 8'h00;
    mem[400] = 8'h00;
    mem[401] = 8'h00;
    mem[402] = 8'h00;
    mem[403] = 8'h00;
    mem[404] = 8'h00;
    mem[405] = 8'h00;
    mem[406] = 8'h00;
    mem[407] = 8'h00;
    mem[408] = 8'h00;
    mem[409] = 8'h00;
    mem[410] = 8'h00;
    mem[411] = 8'h00;
    mem[412] = 8'h00;
    mem[413] = 8'h00;
    mem[414] = 8'h00;
    mem[415] = 8'h00;
    mem[416] = 8'h00;
    mem[417] = 8'h00;
    mem[418] = 8'h00;
    mem[419] = 8'h00;
    mem[420] = 8'h00;
    mem[421] = 8'h00;
    mem[422] = 8'h00;
    mem[423] = 8'h00;
    mem[424] = 8'h00;
    mem[425] = 8'h00;
    mem[426] = 8'h00;
    mem[427] = 8'h00;
    mem[428] = 8'h00;
    mem[429] = 8'h00;
    mem[430] = 8'h00;
    mem[431] = 8'h00;
    mem[432] = 8'h00;
    mem[433] = 8'h00;
    mem[434] = 8'h00;
    mem[435] = 8'h00;
    mem[436] = 8'h00;
    mem[437] = 8'h00;
    mem[438] = 8'h00;
    mem[439] = 8'h00;
    mem[440] = 8'h00;
    mem[441] = 8'h00;
    mem[442] = 8'h00;
    mem[443] = 8'h00;
    mem[444] = 8'h00;
    mem[445] = 8'h00;
    mem[446] = 8'h00;
    mem[447] = 8'h00;
    mem[448] = 8'h00;
    mem[449] = 8'h00;
    mem[450] = 8'h00;
    mem[451] = 8'h00;
    mem[452] = 8'h00;
    mem[453] = 8'h00;
    mem[454] = 8'h00;
    mem[455] = 8'h00;
    mem[456] = 8'h00;
    mem[457] = 8'h00;
    mem[458] = 8'h00;
    mem[459] = 8'h00;
    mem[460] = 8'h00;
    mem[461] = 8'h00;
    mem[462] = 8'h00;
    mem[463] = 8'h00;
    mem[464] = 8'h00;
    mem[465] = 8'h00;
    mem[466] = 8'h00;
    mem[467] = 8'h00;
    mem[468] = 8'h00;
    mem[469] = 8'h00;
    mem[470] = 8'h00;
    mem[471] = 8'h00;
    mem[472] = 8'h00;
    mem[473] = 8'h00;
    mem[474] = 8'h00;
    mem[475] = 8'h00;
    mem[476] = 8'h00;
    mem[477] = 8'h00;
    mem[478] = 8'h00;
    mem[479] = 8'h00;
    mem[480] = 8'h00;
    mem[481] = 8'h00;
    mem[482] = 8'h00;
    mem[483] = 8'h00;
    mem[484] = 8'h00;
    mem[485] = 8'h00;
    mem[486] = 8'h00;
    mem[487] = 8'h00;
    mem[488] = 8'h00;
    mem[489] = 8'h00;
    mem[490] = 8'h00;
    mem[491] = 8'h00;
    mem[492] = 8'h00;
    mem[493] = 8'h00;
    mem[494] = 8'h00;
    mem[495] = 8'h00;
    mem[496] = 8'h00;
    mem[497] = 8'h00;
    mem[498] = 8'h00;
    mem[499] = 8'h00;
    mem[500] = 8'h00;
    mem[501] = 8'h00;
    mem[502] = 8'h00;
    mem[503] = 8'h00;
    mem[504] = 8'h00;
    mem[505] = 8'h00;
    mem[506] = 8'h00;
    mem[507] = 8'h00;
    mem[508] = 8'h00;
    mem[509] = 8'h00;
    mem[510] = 8'h00;
    mem[511] = 8'h00;
  end

  wire [8:0] addr = {y[5:0], x[5:3]};
  assign pixel = mem[addr][x&7];

endmodule

module glyph_512 (
    input wire [5:0] x,
    input wire [5:0] y,
    output wire pixel
);

  reg [7:0] mem[511:0];
  initial begin
    mem[0] = 8'h00;
    mem[1] = 8'h00;
    mem[2] = 8'h00;
    mem[3] = 8'h00;
    mem[4] = 8'h00;
    mem[5] = 8'h00;
    mem[6] = 8'h00;
    mem[7] = 8'h00;
    mem[8] = 8'h00;
    mem[9] = 8'h00;
    mem[10] = 8'h00;
    mem[11] = 8'h00;
    mem[12] = 8'h00;
    mem[13] = 8'h00;
    mem[14] = 8'h00;
    mem[15] = 8'h00;
    mem[16] = 8'h00;
    mem[17] = 8'h00;
    mem[18] = 8'h00;
    mem[19] = 8'h00;
    mem[20] = 8'h00;
    mem[21] = 8'h00;
    mem[22] = 8'h00;
    mem[23] = 8'h00;
    mem[24] = 8'h00;
    mem[25] = 8'h00;
    mem[26] = 8'h00;
    mem[27] = 8'h00;
    mem[28] = 8'h00;
    mem[29] = 8'h00;
    mem[30] = 8'h00;
    mem[31] = 8'h00;
    mem[32] = 8'h00;
    mem[33] = 8'h00;
    mem[34] = 8'h00;
    mem[35] = 8'h00;
    mem[36] = 8'h00;
    mem[37] = 8'h00;
    mem[38] = 8'h00;
    mem[39] = 8'h00;
    mem[40] = 8'h00;
    mem[41] = 8'h00;
    mem[42] = 8'h00;
    mem[43] = 8'h00;
    mem[44] = 8'h00;
    mem[45] = 8'h00;
    mem[46] = 8'h00;
    mem[47] = 8'h00;
    mem[48] = 8'h00;
    mem[49] = 8'h00;
    mem[50] = 8'h00;
    mem[51] = 8'h00;
    mem[52] = 8'h00;
    mem[53] = 8'h00;
    mem[54] = 8'h00;
    mem[55] = 8'h00;
    mem[56] = 8'h00;
    mem[57] = 8'h00;
    mem[58] = 8'h00;
    mem[59] = 8'h00;
    mem[60] = 8'h00;
    mem[61] = 8'h00;
    mem[62] = 8'h00;
    mem[63] = 8'h00;
    mem[64] = 8'h00;
    mem[65] = 8'h00;
    mem[66] = 8'h00;
    mem[67] = 8'h00;
    mem[68] = 8'h00;
    mem[69] = 8'h00;
    mem[70] = 8'h00;
    mem[71] = 8'h00;
    mem[72] = 8'h00;
    mem[73] = 8'h00;
    mem[74] = 8'h00;
    mem[75] = 8'h00;
    mem[76] = 8'h00;
    mem[77] = 8'h00;
    mem[78] = 8'h00;
    mem[79] = 8'h00;
    mem[80] = 8'h00;
    mem[81] = 8'h00;
    mem[82] = 8'h00;
    mem[83] = 8'h00;
    mem[84] = 8'h00;
    mem[85] = 8'h00;
    mem[86] = 8'h00;
    mem[87] = 8'h00;
    mem[88] = 8'h00;
    mem[89] = 8'h00;
    mem[90] = 8'h00;
    mem[91] = 8'h00;
    mem[92] = 8'h00;
    mem[93] = 8'h00;
    mem[94] = 8'h00;
    mem[95] = 8'h00;
    mem[96] = 8'h00;
    mem[97] = 8'h00;
    mem[98] = 8'h00;
    mem[99] = 8'h00;
    mem[100] = 8'h00;
    mem[101] = 8'h00;
    mem[102] = 8'h00;
    mem[103] = 8'h00;
    mem[104] = 8'h00;
    mem[105] = 8'h00;
    mem[106] = 8'h00;
    mem[107] = 8'h00;
    mem[108] = 8'h00;
    mem[109] = 8'h00;
    mem[110] = 8'h00;
    mem[111] = 8'h00;
    mem[112] = 8'h00;
    mem[113] = 8'h00;
    mem[114] = 8'h00;
    mem[115] = 8'h00;
    mem[116] = 8'h00;
    mem[117] = 8'h00;
    mem[118] = 8'h00;
    mem[119] = 8'h00;
    mem[120] = 8'h00;
    mem[121] = 8'h00;
    mem[122] = 8'h00;
    mem[123] = 8'h00;
    mem[124] = 8'h00;
    mem[125] = 8'h00;
    mem[126] = 8'h00;
    mem[127] = 8'h00;
    mem[128] = 8'h00;
    mem[129] = 8'h00;
    mem[130] = 8'h00;
    mem[131] = 8'h00;
    mem[132] = 8'h00;
    mem[133] = 8'h00;
    mem[134] = 8'h00;
    mem[135] = 8'h00;
    mem[136] = 8'h00;
    mem[137] = 8'h00;
    mem[138] = 8'h00;
    mem[139] = 8'h00;
    mem[140] = 8'h00;
    mem[141] = 8'h00;
    mem[142] = 8'h00;
    mem[143] = 8'h00;
    mem[144] = 8'h00;
    mem[145] = 8'h00;
    mem[146] = 8'h00;
    mem[147] = 8'h00;
    mem[148] = 8'h00;
    mem[149] = 8'h00;
    mem[150] = 8'h00;
    mem[151] = 8'h00;
    mem[152] = 8'h00;
    mem[153] = 8'h00;
    mem[154] = 8'h00;
    mem[155] = 8'h00;
    mem[156] = 8'h00;
    mem[157] = 8'h00;
    mem[158] = 8'h00;
    mem[159] = 8'h00;
    mem[160] = 8'hf0;
    mem[161] = 8'hff;
    mem[162] = 8'h03;
    mem[163] = 8'h00;
    mem[164] = 8'h0f;
    mem[165] = 8'h00;
    mem[166] = 8'hfe;
    mem[167] = 8'h03;
    mem[168] = 8'hf0;
    mem[169] = 8'hff;
    mem[170] = 8'h03;
    mem[171] = 8'hc0;
    mem[172] = 8'h0f;
    mem[173] = 8'h80;
    mem[174] = 8'hff;
    mem[175] = 8'h07;
    mem[176] = 8'h70;
    mem[177] = 8'h00;
    mem[178] = 8'h00;
    mem[179] = 8'he0;
    mem[180] = 8'h0f;
    mem[181] = 8'hc0;
    mem[182] = 8'h87;
    mem[183] = 8'h0f;
    mem[184] = 8'h70;
    mem[185] = 8'h00;
    mem[186] = 8'h00;
    mem[187] = 8'hf8;
    mem[188] = 8'h0f;
    mem[189] = 8'hc0;
    mem[190] = 8'h01;
    mem[191] = 8'h0e;
    mem[192] = 8'h70;
    mem[193] = 8'h00;
    mem[194] = 8'h00;
    mem[195] = 8'h7c;
    mem[196] = 8'h0e;
    mem[197] = 8'he0;
    mem[198] = 8'h01;
    mem[199] = 8'h1e;
    mem[200] = 8'h30;
    mem[201] = 8'h00;
    mem[202] = 8'h00;
    mem[203] = 8'h1c;
    mem[204] = 8'h0e;
    mem[205] = 8'he0;
    mem[206] = 8'h00;
    mem[207] = 8'h1e;
    mem[208] = 8'h30;
    mem[209] = 8'h00;
    mem[210] = 8'h00;
    mem[211] = 8'h0c;
    mem[212] = 8'h0e;
    mem[213] = 8'he0;
    mem[214] = 8'h00;
    mem[215] = 8'h1c;
    mem[216] = 8'h38;
    mem[217] = 8'h00;
    mem[218] = 8'h00;
    mem[219] = 8'h00;
    mem[220] = 8'h0e;
    mem[221] = 8'he0;
    mem[222] = 8'h00;
    mem[223] = 8'h1e;
    mem[224] = 8'h38;
    mem[225] = 8'h3f;
    mem[226] = 8'h00;
    mem[227] = 8'h00;
    mem[228] = 8'h0e;
    mem[229] = 8'h00;
    mem[230] = 8'h00;
    mem[231] = 8'h1e;
    mem[232] = 8'hb8;
    mem[233] = 8'hff;
    mem[234] = 8'h00;
    mem[235] = 8'h00;
    mem[236] = 8'h0e;
    mem[237] = 8'h00;
    mem[238] = 8'h00;
    mem[239] = 8'h0e;
    mem[240] = 8'hf8;
    mem[241] = 8'hf3;
    mem[242] = 8'h01;
    mem[243] = 8'h00;
    mem[244] = 8'h0e;
    mem[245] = 8'h00;
    mem[246] = 8'h00;
    mem[247] = 8'h0f;
    mem[248] = 8'hf8;
    mem[249] = 8'hc0;
    mem[250] = 8'h03;
    mem[251] = 8'h00;
    mem[252] = 8'h0e;
    mem[253] = 8'h00;
    mem[254] = 8'h80;
    mem[255] = 8'h07;
    mem[256] = 8'h78;
    mem[257] = 8'h80;
    mem[258] = 8'h07;
    mem[259] = 8'h00;
    mem[260] = 8'h0e;
    mem[261] = 8'h00;
    mem[262] = 8'h80;
    mem[263] = 8'h03;
    mem[264] = 8'h38;
    mem[265] = 8'h80;
    mem[266] = 8'h07;
    mem[267] = 8'h00;
    mem[268] = 8'h0e;
    mem[269] = 8'h00;
    mem[270] = 8'hc0;
    mem[271] = 8'h03;
    mem[272] = 8'h00;
    mem[273] = 8'h00;
    mem[274] = 8'h07;
    mem[275] = 8'h00;
    mem[276] = 8'h0e;
    mem[277] = 8'h00;
    mem[278] = 8'he0;
    mem[279] = 8'h01;
    mem[280] = 8'h00;
    mem[281] = 8'h00;
    mem[282] = 8'h07;
    mem[283] = 8'h00;
    mem[284] = 8'h0e;
    mem[285] = 8'h00;
    mem[286] = 8'hf0;
    mem[287] = 8'h00;
    mem[288] = 8'h00;
    mem[289] = 8'h00;
    mem[290] = 8'h07;
    mem[291] = 8'h00;
    mem[292] = 8'h0e;
    mem[293] = 8'h00;
    mem[294] = 8'h78;
    mem[295] = 8'h00;
    mem[296] = 8'h00;
    mem[297] = 8'h00;
    mem[298] = 8'h07;
    mem[299] = 8'h00;
    mem[300] = 8'h0e;
    mem[301] = 8'h00;
    mem[302] = 8'h3c;
    mem[303] = 8'h00;
    mem[304] = 8'h1c;
    mem[305] = 8'h00;
    mem[306] = 8'h07;
    mem[307] = 8'h00;
    mem[308] = 8'h0e;
    mem[309] = 8'h00;
    mem[310] = 8'h1e;
    mem[311] = 8'h00;
    mem[312] = 8'h3c;
    mem[313] = 8'h00;
    mem[314] = 8'h07;
    mem[315] = 8'h00;
    mem[316] = 8'h0e;
    mem[317] = 8'h00;
    mem[318] = 8'h0f;
    mem[319] = 8'h00;
    mem[320] = 8'h38;
    mem[321] = 8'h80;
    mem[322] = 8'h07;
    mem[323] = 8'h00;
    mem[324] = 8'h0e;
    mem[325] = 8'h80;
    mem[326] = 8'h07;
    mem[327] = 8'h00;
    mem[328] = 8'h78;
    mem[329] = 8'hc0;
    mem[330] = 8'h03;
    mem[331] = 8'h00;
    mem[332] = 8'h0e;
    mem[333] = 8'hc0;
    mem[334] = 8'h03;
    mem[335] = 8'h00;
    mem[336] = 8'hf0;
    mem[337] = 8'he0;
    mem[338] = 8'h01;
    mem[339] = 8'h00;
    mem[340] = 8'h0e;
    mem[341] = 8'he0;
    mem[342] = 8'h01;
    mem[343] = 8'h00;
    mem[344] = 8'he0;
    mem[345] = 8'hff;
    mem[346] = 8'h00;
    mem[347] = 8'h00;
    mem[348] = 8'h0e;
    mem[349] = 8'hf0;
    mem[350] = 8'hff;
    mem[351] = 8'h1f;
    mem[352] = 8'hc0;
    mem[353] = 8'h7f;
    mem[354] = 8'h00;
    mem[355] = 8'h00;
    mem[356] = 8'h0e;
    mem[357] = 8'hf0;
    mem[358] = 8'hff;
    mem[359] = 8'h1f;
    mem[360] = 8'h00;
    mem[361] = 8'h00;
    mem[362] = 8'h00;
    mem[363] = 8'h00;
    mem[364] = 8'h00;
    mem[365] = 8'h00;
    mem[366] = 8'h00;
    mem[367] = 8'h00;
    mem[368] = 8'h00;
    mem[369] = 8'h00;
    mem[370] = 8'h00;
    mem[371] = 8'h00;
    mem[372] = 8'h00;
    mem[373] = 8'h00;
    mem[374] = 8'h00;
    mem[375] = 8'h00;
    mem[376] = 8'h00;
    mem[377] = 8'h00;
    mem[378] = 8'h00;
    mem[379] = 8'h00;
    mem[380] = 8'h00;
    mem[381] = 8'h00;
    mem[382] = 8'h00;
    mem[383] = 8'h00;
    mem[384] = 8'h00;
    mem[385] = 8'h00;
    mem[386] = 8'h00;
    mem[387] = 8'h00;
    mem[388] = 8'h00;
    mem[389] = 8'h00;
    mem[390] = 8'h00;
    mem[391] = 8'h00;
    mem[392] = 8'h00;
    mem[393] = 8'h00;
    mem[394] = 8'h00;
    mem[395] = 8'h00;
    mem[396] = 8'h00;
    mem[397] = 8'h00;
    mem[398] = 8'h00;
    mem[399] = 8'h00;
    mem[400] = 8'h00;
    mem[401] = 8'h00;
    mem[402] = 8'h00;
    mem[403] = 8'h00;
    mem[404] = 8'h00;
    mem[405] = 8'h00;
    mem[406] = 8'h00;
    mem[407] = 8'h00;
    mem[408] = 8'h00;
    mem[409] = 8'h00;
    mem[410] = 8'h00;
    mem[411] = 8'h00;
    mem[412] = 8'h00;
    mem[413] = 8'h00;
    mem[414] = 8'h00;
    mem[415] = 8'h00;
    mem[416] = 8'h00;
    mem[417] = 8'h00;
    mem[418] = 8'h00;
    mem[419] = 8'h00;
    mem[420] = 8'h00;
    mem[421] = 8'h00;
    mem[422] = 8'h00;
    mem[423] = 8'h00;
    mem[424] = 8'h00;
    mem[425] = 8'h00;
    mem[426] = 8'h00;
    mem[427] = 8'h00;
    mem[428] = 8'h00;
    mem[429] = 8'h00;
    mem[430] = 8'h00;
    mem[431] = 8'h00;
    mem[432] = 8'h00;
    mem[433] = 8'h00;
    mem[434] = 8'h00;
    mem[435] = 8'h00;
    mem[436] = 8'h00;
    mem[437] = 8'h00;
    mem[438] = 8'h00;
    mem[439] = 8'h00;
    mem[440] = 8'h00;
    mem[441] = 8'h00;
    mem[442] = 8'h00;
    mem[443] = 8'h00;
    mem[444] = 8'h00;
    mem[445] = 8'h00;
    mem[446] = 8'h00;
    mem[447] = 8'h00;
    mem[448] = 8'h00;
    mem[449] = 8'h00;
    mem[450] = 8'h00;
    mem[451] = 8'h00;
    mem[452] = 8'h00;
    mem[453] = 8'h00;
    mem[454] = 8'h00;
    mem[455] = 8'h00;
    mem[456] = 8'h00;
    mem[457] = 8'h00;
    mem[458] = 8'h00;
    mem[459] = 8'h00;
    mem[460] = 8'h00;
    mem[461] = 8'h00;
    mem[462] = 8'h00;
    mem[463] = 8'h00;
    mem[464] = 8'h00;
    mem[465] = 8'h00;
    mem[466] = 8'h00;
    mem[467] = 8'h00;
    mem[468] = 8'h00;
    mem[469] = 8'h00;
    mem[470] = 8'h00;
    mem[471] = 8'h00;
    mem[472] = 8'h00;
    mem[473] = 8'h00;
    mem[474] = 8'h00;
    mem[475] = 8'h00;
    mem[476] = 8'h00;
    mem[477] = 8'h00;
    mem[478] = 8'h00;
    mem[479] = 8'h00;
    mem[480] = 8'h00;
    mem[481] = 8'h00;
    mem[482] = 8'h00;
    mem[483] = 8'h00;
    mem[484] = 8'h00;
    mem[485] = 8'h00;
    mem[486] = 8'h00;
    mem[487] = 8'h00;
    mem[488] = 8'h00;
    mem[489] = 8'h00;
    mem[490] = 8'h00;
    mem[491] = 8'h00;
    mem[492] = 8'h00;
    mem[493] = 8'h00;
    mem[494] = 8'h00;
    mem[495] = 8'h00;
    mem[496] = 8'h00;
    mem[497] = 8'h00;
    mem[498] = 8'h00;
    mem[499] = 8'h00;
    mem[500] = 8'h00;
    mem[501] = 8'h00;
    mem[502] = 8'h00;
    mem[503] = 8'h00;
    mem[504] = 8'h00;
    mem[505] = 8'h00;
    mem[506] = 8'h00;
    mem[507] = 8'h00;
    mem[508] = 8'h00;
    mem[509] = 8'h00;
    mem[510] = 8'h00;
    mem[511] = 8'h00;
  end

  wire [8:0] addr = {y[5:0], x[5:3]};
  assign pixel = mem[addr][x&7];

endmodule

module glyph_1024 (
    input wire [5:0] x,
    input wire [5:0] y,
    output wire pixel
);

  reg [7:0] mem[511:0];
  initial begin
    mem[0] = 8'h00;
    mem[1] = 8'h00;
    mem[2] = 8'h00;
    mem[3] = 8'h00;
    mem[4] = 8'h00;
    mem[5] = 8'h00;
    mem[6] = 8'h00;
    mem[7] = 8'h00;
    mem[8] = 8'h00;
    mem[9] = 8'h00;
    mem[10] = 8'h00;
    mem[11] = 8'h00;
    mem[12] = 8'h00;
    mem[13] = 8'h00;
    mem[14] = 8'h00;
    mem[15] = 8'h00;
    mem[16] = 8'h00;
    mem[17] = 8'h00;
    mem[18] = 8'h00;
    mem[19] = 8'h00;
    mem[20] = 8'h00;
    mem[21] = 8'h00;
    mem[22] = 8'h00;
    mem[23] = 8'h00;
    mem[24] = 8'h00;
    mem[25] = 8'h00;
    mem[26] = 8'h00;
    mem[27] = 8'h00;
    mem[28] = 8'h00;
    mem[29] = 8'h00;
    mem[30] = 8'h00;
    mem[31] = 8'h00;
    mem[32] = 8'h00;
    mem[33] = 8'h00;
    mem[34] = 8'h00;
    mem[35] = 8'h00;
    mem[36] = 8'h00;
    mem[37] = 8'h00;
    mem[38] = 8'h00;
    mem[39] = 8'h00;
    mem[40] = 8'h00;
    mem[41] = 8'h00;
    mem[42] = 8'h00;
    mem[43] = 8'h00;
    mem[44] = 8'h00;
    mem[45] = 8'h00;
    mem[46] = 8'h00;
    mem[47] = 8'h00;
    mem[48] = 8'h00;
    mem[49] = 8'h00;
    mem[50] = 8'h00;
    mem[51] = 8'h00;
    mem[52] = 8'h00;
    mem[53] = 8'h00;
    mem[54] = 8'h00;
    mem[55] = 8'h00;
    mem[56] = 8'h00;
    mem[57] = 8'h00;
    mem[58] = 8'h00;
    mem[59] = 8'h00;
    mem[60] = 8'h00;
    mem[61] = 8'h00;
    mem[62] = 8'h00;
    mem[63] = 8'h00;
    mem[64] = 8'h00;
    mem[65] = 8'h00;
    mem[66] = 8'h00;
    mem[67] = 8'h00;
    mem[68] = 8'h00;
    mem[69] = 8'h00;
    mem[70] = 8'h00;
    mem[71] = 8'h00;
    mem[72] = 8'h00;
    mem[73] = 8'h00;
    mem[74] = 8'h00;
    mem[75] = 8'h00;
    mem[76] = 8'h00;
    mem[77] = 8'h00;
    mem[78] = 8'h00;
    mem[79] = 8'h00;
    mem[80] = 8'h00;
    mem[81] = 8'h00;
    mem[82] = 8'h00;
    mem[83] = 8'h00;
    mem[84] = 8'h00;
    mem[85] = 8'h00;
    mem[86] = 8'h00;
    mem[87] = 8'h00;
    mem[88] = 8'h00;
    mem[89] = 8'h00;
    mem[90] = 8'h00;
    mem[91] = 8'h00;
    mem[92] = 8'h00;
    mem[93] = 8'h00;
    mem[94] = 8'h00;
    mem[95] = 8'h00;
    mem[96] = 8'h00;
    mem[97] = 8'h00;
    mem[98] = 8'h00;
    mem[99] = 8'h00;
    mem[100] = 8'h00;
    mem[101] = 8'h00;
    mem[102] = 8'h00;
    mem[103] = 8'h00;
    mem[104] = 8'h00;
    mem[105] = 8'h00;
    mem[106] = 8'h00;
    mem[107] = 8'h00;
    mem[108] = 8'h00;
    mem[109] = 8'h00;
    mem[110] = 8'h00;
    mem[111] = 8'h00;
    mem[112] = 8'h00;
    mem[113] = 8'h00;
    mem[114] = 8'h00;
    mem[115] = 8'h00;
    mem[116] = 8'h00;
    mem[117] = 8'h00;
    mem[118] = 8'h00;
    mem[119] = 8'h00;
    mem[120] = 8'h00;
    mem[121] = 8'h00;
    mem[122] = 8'h00;
    mem[123] = 8'h00;
    mem[124] = 8'h00;
    mem[125] = 8'h00;
    mem[126] = 8'h00;
    mem[127] = 8'h00;
    mem[128] = 8'h00;
    mem[129] = 8'h00;
    mem[130] = 8'h00;
    mem[131] = 8'h00;
    mem[132] = 8'h00;
    mem[133] = 8'h00;
    mem[134] = 8'h00;
    mem[135] = 8'h00;
    mem[136] = 8'h00;
    mem[137] = 8'h00;
    mem[138] = 8'h00;
    mem[139] = 8'h00;
    mem[140] = 8'h00;
    mem[141] = 8'h00;
    mem[142] = 8'h00;
    mem[143] = 8'h00;
    mem[144] = 8'h00;
    mem[145] = 8'h00;
    mem[146] = 8'h00;
    mem[147] = 8'h00;
    mem[148] = 8'h00;
    mem[149] = 8'h00;
    mem[150] = 8'h00;
    mem[151] = 8'h00;
    mem[152] = 8'h00;
    mem[153] = 8'h00;
    mem[154] = 8'h00;
    mem[155] = 8'h00;
    mem[156] = 8'h00;
    mem[157] = 8'h00;
    mem[158] = 8'h00;
    mem[159] = 8'h00;
    mem[160] = 8'h00;
    mem[161] = 8'h00;
    mem[162] = 8'h00;
    mem[163] = 8'h00;
    mem[164] = 8'h00;
    mem[165] = 8'h00;
    mem[166] = 8'h00;
    mem[167] = 8'h00;
    mem[168] = 8'h00;
    mem[169] = 8'h00;
    mem[170] = 8'h00;
    mem[171] = 8'h00;
    mem[172] = 8'h00;
    mem[173] = 8'h00;
    mem[174] = 8'h00;
    mem[175] = 8'h00;
    mem[176] = 8'h00;
    mem[177] = 8'h00;
    mem[178] = 8'h00;
    mem[179] = 8'h00;
    mem[180] = 8'h00;
    mem[181] = 8'h00;
    mem[182] = 8'h00;
    mem[183] = 8'h00;
    mem[184] = 8'h00;
    mem[185] = 8'h00;
    mem[186] = 8'h00;
    mem[187] = 8'h00;
    mem[188] = 8'h00;
    mem[189] = 8'h00;
    mem[190] = 8'h00;
    mem[191] = 8'h00;
    mem[192] = 8'h00;
    mem[193] = 8'h0f;
    mem[194] = 8'he0;
    mem[195] = 8'h07;
    mem[196] = 8'hc0;
    mem[197] = 8'h0f;
    mem[198] = 8'h00;
    mem[199] = 8'h1c;
    mem[200] = 8'hc0;
    mem[201] = 8'h0f;
    mem[202] = 8'hf0;
    mem[203] = 8'h0f;
    mem[204] = 8'he0;
    mem[205] = 8'h1f;
    mem[206] = 8'h00;
    mem[207] = 8'h1e;
    mem[208] = 8'he0;
    mem[209] = 8'h0f;
    mem[210] = 8'h38;
    mem[211] = 8'h1c;
    mem[212] = 8'h70;
    mem[213] = 8'h38;
    mem[214] = 8'h00;
    mem[215] = 8'h1e;
    mem[216] = 8'h70;
    mem[217] = 8'h0e;
    mem[218] = 8'h1c;
    mem[219] = 8'h38;
    mem[220] = 8'h38;
    mem[221] = 8'h70;
    mem[222] = 8'h00;
    mem[223] = 8'h1f;
    mem[224] = 8'h18;
    mem[225] = 8'h0e;
    mem[226] = 8'h0c;
    mem[227] = 8'h30;
    mem[228] = 8'h18;
    mem[229] = 8'h70;
    mem[230] = 8'h80;
    mem[231] = 8'h1f;
    mem[232] = 8'h00;
    mem[233] = 8'h0e;
    mem[234] = 8'h0e;
    mem[235] = 8'h70;
    mem[236] = 8'h18;
    mem[237] = 8'h70;
    mem[238] = 8'hc0;
    mem[239] = 8'h1d;
    mem[240] = 8'h00;
    mem[241] = 8'h0e;
    mem[242] = 8'h0e;
    mem[243] = 8'h70;
    mem[244] = 8'h00;
    mem[245] = 8'h70;
    mem[246] = 8'hc0;
    mem[247] = 8'h1c;
    mem[248] = 8'h00;
    mem[249] = 8'h0e;
    mem[250] = 8'h0e;
    mem[251] = 8'h70;
    mem[252] = 8'h00;
    mem[253] = 8'h30;
    mem[254] = 8'h60;
    mem[255] = 8'h1c;
    mem[256] = 8'h00;
    mem[257] = 8'h0e;
    mem[258] = 8'h0e;
    mem[259] = 8'h70;
    mem[260] = 8'h00;
    mem[261] = 8'h38;
    mem[262] = 8'h70;
    mem[263] = 8'h1c;
    mem[264] = 8'h00;
    mem[265] = 8'h0e;
    mem[266] = 8'h0e;
    mem[267] = 8'h70;
    mem[268] = 8'h00;
    mem[269] = 8'h1c;
    mem[270] = 8'h38;
    mem[271] = 8'h1c;
    mem[272] = 8'h00;
    mem[273] = 8'h0e;
    mem[274] = 8'h0e;
    mem[275] = 8'h70;
    mem[276] = 8'h00;
    mem[277] = 8'h0e;
    mem[278] = 8'h18;
    mem[279] = 8'h1c;
    mem[280] = 8'h00;
    mem[281] = 8'h0e;
    mem[282] = 8'h0e;
    mem[283] = 8'h70;
    mem[284] = 8'h00;
    mem[285] = 8'h07;
    mem[286] = 8'h0c;
    mem[287] = 8'h1c;
    mem[288] = 8'h00;
    mem[289] = 8'h0e;
    mem[290] = 8'h0e;
    mem[291] = 8'h70;
    mem[292] = 8'h80;
    mem[293] = 8'h03;
    mem[294] = 8'hfe;
    mem[295] = 8'h7f;
    mem[296] = 8'h00;
    mem[297] = 8'h0e;
    mem[298] = 8'h0e;
    mem[299] = 8'h70;
    mem[300] = 8'hc0;
    mem[301] = 8'h01;
    mem[302] = 8'hfe;
    mem[303] = 8'h7f;
    mem[304] = 8'h00;
    mem[305] = 8'h0e;
    mem[306] = 8'h0c;
    mem[307] = 8'h30;
    mem[308] = 8'he0;
    mem[309] = 8'h00;
    mem[310] = 8'h00;
    mem[311] = 8'h1c;
    mem[312] = 8'h00;
    mem[313] = 8'h0e;
    mem[314] = 8'h1c;
    mem[315] = 8'h38;
    mem[316] = 8'h70;
    mem[317] = 8'h00;
    mem[318] = 8'h00;
    mem[319] = 8'h1c;
    mem[320] = 8'h00;
    mem[321] = 8'h0e;
    mem[322] = 8'h38;
    mem[323] = 8'h1c;
    mem[324] = 8'h38;
    mem[325] = 8'h00;
    mem[326] = 8'h00;
    mem[327] = 8'h1c;
    mem[328] = 8'h00;
    mem[329] = 8'h0e;
    mem[330] = 8'hf0;
    mem[331] = 8'h0f;
    mem[332] = 8'hfc;
    mem[333] = 8'h7f;
    mem[334] = 8'h00;
    mem[335] = 8'h1c;
    mem[336] = 8'h00;
    mem[337] = 8'h0e;
    mem[338] = 8'he0;
    mem[339] = 8'h07;
    mem[340] = 8'hfc;
    mem[341] = 8'h7f;
    mem[342] = 8'h00;
    mem[343] = 8'h1c;
    mem[344] = 8'h00;
    mem[345] = 8'h00;
    mem[346] = 8'h00;
    mem[347] = 8'h00;
    mem[348] = 8'h00;
    mem[349] = 8'h00;
    mem[350] = 8'h00;
    mem[351] = 8'h00;
    mem[352] = 8'h00;
    mem[353] = 8'h00;
    mem[354] = 8'h00;
    mem[355] = 8'h00;
    mem[356] = 8'h00;
    mem[357] = 8'h00;
    mem[358] = 8'h00;
    mem[359] = 8'h00;
    mem[360] = 8'h00;
    mem[361] = 8'h00;
    mem[362] = 8'h00;
    mem[363] = 8'h00;
    mem[364] = 8'h00;
    mem[365] = 8'h00;
    mem[366] = 8'h00;
    mem[367] = 8'h00;
    mem[368] = 8'h00;
    mem[369] = 8'h00;
    mem[370] = 8'h00;
    mem[371] = 8'h00;
    mem[372] = 8'h00;
    mem[373] = 8'h00;
    mem[374] = 8'h00;
    mem[375] = 8'h00;
    mem[376] = 8'h00;
    mem[377] = 8'h00;
    mem[378] = 8'h00;
    mem[379] = 8'h00;
    mem[380] = 8'h00;
    mem[381] = 8'h00;
    mem[382] = 8'h00;
    mem[383] = 8'h00;
    mem[384] = 8'h00;
    mem[385] = 8'h00;
    mem[386] = 8'h00;
    mem[387] = 8'h00;
    mem[388] = 8'h00;
    mem[389] = 8'h00;
    mem[390] = 8'h00;
    mem[391] = 8'h00;
    mem[392] = 8'h00;
    mem[393] = 8'h00;
    mem[394] = 8'h00;
    mem[395] = 8'h00;
    mem[396] = 8'h00;
    mem[397] = 8'h00;
    mem[398] = 8'h00;
    mem[399] = 8'h00;
    mem[400] = 8'h00;
    mem[401] = 8'h00;
    mem[402] = 8'h00;
    mem[403] = 8'h00;
    mem[404] = 8'h00;
    mem[405] = 8'h00;
    mem[406] = 8'h00;
    mem[407] = 8'h00;
    mem[408] = 8'h00;
    mem[409] = 8'h00;
    mem[410] = 8'h00;
    mem[411] = 8'h00;
    mem[412] = 8'h00;
    mem[413] = 8'h00;
    mem[414] = 8'h00;
    mem[415] = 8'h00;
    mem[416] = 8'h00;
    mem[417] = 8'h00;
    mem[418] = 8'h00;
    mem[419] = 8'h00;
    mem[420] = 8'h00;
    mem[421] = 8'h00;
    mem[422] = 8'h00;
    mem[423] = 8'h00;
    mem[424] = 8'h00;
    mem[425] = 8'h00;
    mem[426] = 8'h00;
    mem[427] = 8'h00;
    mem[428] = 8'h00;
    mem[429] = 8'h00;
    mem[430] = 8'h00;
    mem[431] = 8'h00;
    mem[432] = 8'h00;
    mem[433] = 8'h00;
    mem[434] = 8'h00;
    mem[435] = 8'h00;
    mem[436] = 8'h00;
    mem[437] = 8'h00;
    mem[438] = 8'h00;
    mem[439] = 8'h00;
    mem[440] = 8'h00;
    mem[441] = 8'h00;
    mem[442] = 8'h00;
    mem[443] = 8'h00;
    mem[444] = 8'h00;
    mem[445] = 8'h00;
    mem[446] = 8'h00;
    mem[447] = 8'h00;
    mem[448] = 8'h00;
    mem[449] = 8'h00;
    mem[450] = 8'h00;
    mem[451] = 8'h00;
    mem[452] = 8'h00;
    mem[453] = 8'h00;
    mem[454] = 8'h00;
    mem[455] = 8'h00;
    mem[456] = 8'h00;
    mem[457] = 8'h00;
    mem[458] = 8'h00;
    mem[459] = 8'h00;
    mem[460] = 8'h00;
    mem[461] = 8'h00;
    mem[462] = 8'h00;
    mem[463] = 8'h00;
    mem[464] = 8'h00;
    mem[465] = 8'h00;
    mem[466] = 8'h00;
    mem[467] = 8'h00;
    mem[468] = 8'h00;
    mem[469] = 8'h00;
    mem[470] = 8'h00;
    mem[471] = 8'h00;
    mem[472] = 8'h00;
    mem[473] = 8'h00;
    mem[474] = 8'h00;
    mem[475] = 8'h00;
    mem[476] = 8'h00;
    mem[477] = 8'h00;
    mem[478] = 8'h00;
    mem[479] = 8'h00;
    mem[480] = 8'h00;
    mem[481] = 8'h00;
    mem[482] = 8'h00;
    mem[483] = 8'h00;
    mem[484] = 8'h00;
    mem[485] = 8'h00;
    mem[486] = 8'h00;
    mem[487] = 8'h00;
    mem[488] = 8'h00;
    mem[489] = 8'h00;
    mem[490] = 8'h00;
    mem[491] = 8'h00;
    mem[492] = 8'h00;
    mem[493] = 8'h00;
    mem[494] = 8'h00;
    mem[495] = 8'h00;
    mem[496] = 8'h00;
    mem[497] = 8'h00;
    mem[498] = 8'h00;
    mem[499] = 8'h00;
    mem[500] = 8'h00;
    mem[501] = 8'h00;
    mem[502] = 8'h00;
    mem[503] = 8'h00;
    mem[504] = 8'h00;
    mem[505] = 8'h00;
    mem[506] = 8'h00;
    mem[507] = 8'h00;
    mem[508] = 8'h00;
    mem[509] = 8'h00;
    mem[510] = 8'h00;
    mem[511] = 8'h00;
  end

  wire [8:0] addr = {y[5:0], x[5:3]};
  assign pixel = mem[addr][x&7];

endmodule

module glyph_2048 (
    input wire [5:0] x,
    input wire [5:0] y,
    output wire pixel
);

  reg [7:0] mem[511:0];
  initial begin
    mem[0] = 8'h00;
    mem[1] = 8'h00;
    mem[2] = 8'h00;
    mem[3] = 8'h00;
    mem[4] = 8'h00;
    mem[5] = 8'h00;
    mem[6] = 8'h00;
    mem[7] = 8'h00;
    mem[8] = 8'h00;
    mem[9] = 8'h00;
    mem[10] = 8'h00;
    mem[11] = 8'h00;
    mem[12] = 8'h00;
    mem[13] = 8'h00;
    mem[14] = 8'h00;
    mem[15] = 8'h00;
    mem[16] = 8'h00;
    mem[17] = 8'h00;
    mem[18] = 8'h00;
    mem[19] = 8'h00;
    mem[20] = 8'h00;
    mem[21] = 8'h00;
    mem[22] = 8'h00;
    mem[23] = 8'h00;
    mem[24] = 8'h00;
    mem[25] = 8'h00;
    mem[26] = 8'h00;
    mem[27] = 8'h00;
    mem[28] = 8'h00;
    mem[29] = 8'h00;
    mem[30] = 8'h00;
    mem[31] = 8'h00;
    mem[32] = 8'h00;
    mem[33] = 8'h00;
    mem[34] = 8'h00;
    mem[35] = 8'h00;
    mem[36] = 8'h00;
    mem[37] = 8'h00;
    mem[38] = 8'h00;
    mem[39] = 8'h00;
    mem[40] = 8'h00;
    mem[41] = 8'h00;
    mem[42] = 8'h00;
    mem[43] = 8'h00;
    mem[44] = 8'h00;
    mem[45] = 8'h00;
    mem[46] = 8'h00;
    mem[47] = 8'h00;
    mem[48] = 8'h00;
    mem[49] = 8'h00;
    mem[50] = 8'h00;
    mem[51] = 8'h00;
    mem[52] = 8'h00;
    mem[53] = 8'h00;
    mem[54] = 8'h00;
    mem[55] = 8'h00;
    mem[56] = 8'h00;
    mem[57] = 8'h00;
    mem[58] = 8'h00;
    mem[59] = 8'h00;
    mem[60] = 8'h00;
    mem[61] = 8'h00;
    mem[62] = 8'h00;
    mem[63] = 8'h00;
    mem[64] = 8'h00;
    mem[65] = 8'h00;
    mem[66] = 8'h00;
    mem[67] = 8'h00;
    mem[68] = 8'h00;
    mem[69] = 8'h00;
    mem[70] = 8'h00;
    mem[71] = 8'h00;
    mem[72] = 8'h00;
    mem[73] = 8'h00;
    mem[74] = 8'h00;
    mem[75] = 8'h00;
    mem[76] = 8'h00;
    mem[77] = 8'h00;
    mem[78] = 8'h00;
    mem[79] = 8'h00;
    mem[80] = 8'h00;
    mem[81] = 8'h00;
    mem[82] = 8'h00;
    mem[83] = 8'h00;
    mem[84] = 8'h00;
    mem[85] = 8'h00;
    mem[86] = 8'h00;
    mem[87] = 8'h00;
    mem[88] = 8'h00;
    mem[89] = 8'h00;
    mem[90] = 8'h00;
    mem[91] = 8'h00;
    mem[92] = 8'h00;
    mem[93] = 8'h00;
    mem[94] = 8'h00;
    mem[95] = 8'h00;
    mem[96] = 8'h00;
    mem[97] = 8'h00;
    mem[98] = 8'h00;
    mem[99] = 8'h00;
    mem[100] = 8'h00;
    mem[101] = 8'h00;
    mem[102] = 8'h00;
    mem[103] = 8'h00;
    mem[104] = 8'h00;
    mem[105] = 8'h00;
    mem[106] = 8'h00;
    mem[107] = 8'h00;
    mem[108] = 8'h00;
    mem[109] = 8'h00;
    mem[110] = 8'h00;
    mem[111] = 8'h00;
    mem[112] = 8'h00;
    mem[113] = 8'h00;
    mem[114] = 8'h00;
    mem[115] = 8'h00;
    mem[116] = 8'h00;
    mem[117] = 8'h00;
    mem[118] = 8'h00;
    mem[119] = 8'h00;
    mem[120] = 8'h00;
    mem[121] = 8'h00;
    mem[122] = 8'h00;
    mem[123] = 8'h00;
    mem[124] = 8'h00;
    mem[125] = 8'h00;
    mem[126] = 8'h00;
    mem[127] = 8'h00;
    mem[128] = 8'h00;
    mem[129] = 8'h00;
    mem[130] = 8'h00;
    mem[131] = 8'h00;
    mem[132] = 8'h00;
    mem[133] = 8'h00;
    mem[134] = 8'h00;
    mem[135] = 8'h00;
    mem[136] = 8'h00;
    mem[137] = 8'h00;
    mem[138] = 8'h00;
    mem[139] = 8'h00;
    mem[140] = 8'h00;
    mem[141] = 8'h00;
    mem[142] = 8'h00;
    mem[143] = 8'h00;
    mem[144] = 8'h00;
    mem[145] = 8'h00;
    mem[146] = 8'h00;
    mem[147] = 8'h00;
    mem[148] = 8'h00;
    mem[149] = 8'h00;
    mem[150] = 8'h00;
    mem[151] = 8'h00;
    mem[152] = 8'h00;
    mem[153] = 8'h00;
    mem[154] = 8'h00;
    mem[155] = 8'h00;
    mem[156] = 8'h00;
    mem[157] = 8'h00;
    mem[158] = 8'h00;
    mem[159] = 8'h00;
    mem[160] = 8'h00;
    mem[161] = 8'h00;
    mem[162] = 8'h00;
    mem[163] = 8'h00;
    mem[164] = 8'h00;
    mem[165] = 8'h00;
    mem[166] = 8'h00;
    mem[167] = 8'h00;
    mem[168] = 8'h00;
    mem[169] = 8'h00;
    mem[170] = 8'h00;
    mem[171] = 8'h00;
    mem[172] = 8'h00;
    mem[173] = 8'h00;
    mem[174] = 8'h00;
    mem[175] = 8'h00;
    mem[176] = 8'h00;
    mem[177] = 8'h00;
    mem[178] = 8'h00;
    mem[179] = 8'h00;
    mem[180] = 8'h00;
    mem[181] = 8'h00;
    mem[182] = 8'h00;
    mem[183] = 8'h00;
    mem[184] = 8'h00;
    mem[185] = 8'h00;
    mem[186] = 8'h00;
    mem[187] = 8'h00;
    mem[188] = 8'h00;
    mem[189] = 8'h00;
    mem[190] = 8'h00;
    mem[191] = 8'h00;
    mem[192] = 8'hc0;
    mem[193] = 8'h0f;
    mem[194] = 8'he0;
    mem[195] = 8'h07;
    mem[196] = 8'h00;
    mem[197] = 8'h1c;
    mem[198] = 8'he0;
    mem[199] = 8'h07;
    mem[200] = 8'he0;
    mem[201] = 8'h1f;
    mem[202] = 8'hf0;
    mem[203] = 8'h0f;
    mem[204] = 8'h00;
    mem[205] = 8'h1e;
    mem[206] = 8'hf8;
    mem[207] = 8'h0f;
    mem[208] = 8'h70;
    mem[209] = 8'h38;
    mem[210] = 8'h38;
    mem[211] = 8'h1c;
    mem[212] = 8'h00;
    mem[213] = 8'h1e;
    mem[214] = 8'h38;
    mem[215] = 8'h1c;
    mem[216] = 8'h38;
    mem[217] = 8'h70;
    mem[218] = 8'h1c;
    mem[219] = 8'h38;
    mem[220] = 8'h00;
    mem[221] = 8'h1f;
    mem[222] = 8'h1c;
    mem[223] = 8'h38;
    mem[224] = 8'h18;
    mem[225] = 8'h70;
    mem[226] = 8'h0c;
    mem[227] = 8'h30;
    mem[228] = 8'h80;
    mem[229] = 8'h1f;
    mem[230] = 8'h1c;
    mem[231] = 8'h38;
    mem[232] = 8'h18;
    mem[233] = 8'h70;
    mem[234] = 8'h0e;
    mem[235] = 8'h70;
    mem[236] = 8'hc0;
    mem[237] = 8'h1d;
    mem[238] = 8'h1c;
    mem[239] = 8'h38;
    mem[240] = 8'h00;
    mem[241] = 8'h70;
    mem[242] = 8'h0e;
    mem[243] = 8'h70;
    mem[244] = 8'hc0;
    mem[245] = 8'h1c;
    mem[246] = 8'h1c;
    mem[247] = 8'h38;
    mem[248] = 8'h00;
    mem[249] = 8'h30;
    mem[250] = 8'h0e;
    mem[251] = 8'h70;
    mem[252] = 8'h60;
    mem[253] = 8'h1c;
    mem[254] = 8'h38;
    mem[255] = 8'h1c;
    mem[256] = 8'h00;
    mem[257] = 8'h38;
    mem[258] = 8'h0e;
    mem[259] = 8'h70;
    mem[260] = 8'h70;
    mem[261] = 8'h1c;
    mem[262] = 8'hf0;
    mem[263] = 8'h0f;
    mem[264] = 8'h00;
    mem[265] = 8'h1c;
    mem[266] = 8'h0e;
    mem[267] = 8'h70;
    mem[268] = 8'h38;
    mem[269] = 8'h1c;
    mem[270] = 8'hf8;
    mem[271] = 8'h0f;
    mem[272] = 8'h00;
    mem[273] = 8'h0e;
    mem[274] = 8'h0e;
    mem[275] = 8'h70;
    mem[276] = 8'h18;
    mem[277] = 8'h1c;
    mem[278] = 8'h1c;
    mem[279] = 8'h1c;
    mem[280] = 8'h00;
    mem[281] = 8'h07;
    mem[282] = 8'h0e;
    mem[283] = 8'h70;
    mem[284] = 8'h0c;
    mem[285] = 8'h1c;
    mem[286] = 8'h0e;
    mem[287] = 8'h38;
    mem[288] = 8'h80;
    mem[289] = 8'h03;
    mem[290] = 8'h0e;
    mem[291] = 8'h70;
    mem[292] = 8'hfe;
    mem[293] = 8'h7f;
    mem[294] = 8'h0e;
    mem[295] = 8'h30;
    mem[296] = 8'hc0;
    mem[297] = 8'h01;
    mem[298] = 8'h0e;
    mem[299] = 8'h70;
    mem[300] = 8'hfe;
    mem[301] = 8'h7f;
    mem[302] = 8'h0e;
    mem[303] = 8'h70;
    mem[304] = 8'he0;
    mem[305] = 8'h00;
    mem[306] = 8'h0c;
    mem[307] = 8'h30;
    mem[308] = 8'h00;
    mem[309] = 8'h1c;
    mem[310] = 8'h0e;
    mem[311] = 8'h70;
    mem[312] = 8'h70;
    mem[313] = 8'h00;
    mem[314] = 8'h1c;
    mem[315] = 8'h38;
    mem[316] = 8'h00;
    mem[317] = 8'h1c;
    mem[318] = 8'h0e;
    mem[319] = 8'h38;
    mem[320] = 8'h38;
    mem[321] = 8'h00;
    mem[322] = 8'h38;
    mem[323] = 8'h1c;
    mem[324] = 8'h00;
    mem[325] = 8'h1c;
    mem[326] = 8'h1c;
    mem[327] = 8'h3c;
    mem[328] = 8'hfc;
    mem[329] = 8'h7f;
    mem[330] = 8'hf0;
    mem[331] = 8'h0f;
    mem[332] = 8'h00;
    mem[333] = 8'h1c;
    mem[334] = 8'hf8;
    mem[335] = 8'h1f;
    mem[336] = 8'hfc;
    mem[337] = 8'h7f;
    mem[338] = 8'he0;
    mem[339] = 8'h07;
    mem[340] = 8'h00;
    mem[341] = 8'h1c;
    mem[342] = 8'he0;
    mem[343] = 8'h07;
    mem[344] = 8'h00;
    mem[345] = 8'h00;
    mem[346] = 8'h00;
    mem[347] = 8'h00;
    mem[348] = 8'h00;
    mem[349] = 8'h00;
    mem[350] = 8'h00;
    mem[351] = 8'h00;
    mem[352] = 8'h00;
    mem[353] = 8'h00;
    mem[354] = 8'h00;
    mem[355] = 8'h00;
    mem[356] = 8'h00;
    mem[357] = 8'h00;
    mem[358] = 8'h00;
    mem[359] = 8'h00;
    mem[360] = 8'h00;
    mem[361] = 8'h00;
    mem[362] = 8'h00;
    mem[363] = 8'h00;
    mem[364] = 8'h00;
    mem[365] = 8'h00;
    mem[366] = 8'h00;
    mem[367] = 8'h00;
    mem[368] = 8'h00;
    mem[369] = 8'h00;
    mem[370] = 8'h00;
    mem[371] = 8'h00;
    mem[372] = 8'h00;
    mem[373] = 8'h00;
    mem[374] = 8'h00;
    mem[375] = 8'h00;
    mem[376] = 8'h00;
    mem[377] = 8'h00;
    mem[378] = 8'h00;
    mem[379] = 8'h00;
    mem[380] = 8'h00;
    mem[381] = 8'h00;
    mem[382] = 8'h00;
    mem[383] = 8'h00;
    mem[384] = 8'h00;
    mem[385] = 8'h00;
    mem[386] = 8'h00;
    mem[387] = 8'h00;
    mem[388] = 8'h00;
    mem[389] = 8'h00;
    mem[390] = 8'h00;
    mem[391] = 8'h00;
    mem[392] = 8'h00;
    mem[393] = 8'h00;
    mem[394] = 8'h00;
    mem[395] = 8'h00;
    mem[396] = 8'h00;
    mem[397] = 8'h00;
    mem[398] = 8'h00;
    mem[399] = 8'h00;
    mem[400] = 8'h00;
    mem[401] = 8'h00;
    mem[402] = 8'h00;
    mem[403] = 8'h00;
    mem[404] = 8'h00;
    mem[405] = 8'h00;
    mem[406] = 8'h00;
    mem[407] = 8'h00;
    mem[408] = 8'h00;
    mem[409] = 8'h00;
    mem[410] = 8'h00;
    mem[411] = 8'h00;
    mem[412] = 8'h00;
    mem[413] = 8'h00;
    mem[414] = 8'h00;
    mem[415] = 8'h00;
    mem[416] = 8'h00;
    mem[417] = 8'h00;
    mem[418] = 8'h00;
    mem[419] = 8'h00;
    mem[420] = 8'h00;
    mem[421] = 8'h00;
    mem[422] = 8'h00;
    mem[423] = 8'h00;
    mem[424] = 8'h00;
    mem[425] = 8'h00;
    mem[426] = 8'h00;
    mem[427] = 8'h00;
    mem[428] = 8'h00;
    mem[429] = 8'h00;
    mem[430] = 8'h00;
    mem[431] = 8'h00;
    mem[432] = 8'h00;
    mem[433] = 8'h00;
    mem[434] = 8'h00;
    mem[435] = 8'h00;
    mem[436] = 8'h00;
    mem[437] = 8'h00;
    mem[438] = 8'h00;
    mem[439] = 8'h00;
    mem[440] = 8'h00;
    mem[441] = 8'h00;
    mem[442] = 8'h00;
    mem[443] = 8'h00;
    mem[444] = 8'h00;
    mem[445] = 8'h00;
    mem[446] = 8'h00;
    mem[447] = 8'h00;
    mem[448] = 8'h00;
    mem[449] = 8'h00;
    mem[450] = 8'h00;
    mem[451] = 8'h00;
    mem[452] = 8'h00;
    mem[453] = 8'h00;
    mem[454] = 8'h00;
    mem[455] = 8'h00;
    mem[456] = 8'h00;
    mem[457] = 8'h00;
    mem[458] = 8'h00;
    mem[459] = 8'h00;
    mem[460] = 8'h00;
    mem[461] = 8'h00;
    mem[462] = 8'h00;
    mem[463] = 8'h00;
    mem[464] = 8'h00;
    mem[465] = 8'h00;
    mem[466] = 8'h00;
    mem[467] = 8'h00;
    mem[468] = 8'h00;
    mem[469] = 8'h00;
    mem[470] = 8'h00;
    mem[471] = 8'h00;
    mem[472] = 8'h00;
    mem[473] = 8'h00;
    mem[474] = 8'h00;
    mem[475] = 8'h00;
    mem[476] = 8'h00;
    mem[477] = 8'h00;
    mem[478] = 8'h00;
    mem[479] = 8'h00;
    mem[480] = 8'h00;
    mem[481] = 8'h00;
    mem[482] = 8'h00;
    mem[483] = 8'h00;
    mem[484] = 8'h00;
    mem[485] = 8'h00;
    mem[486] = 8'h00;
    mem[487] = 8'h00;
    mem[488] = 8'h00;
    mem[489] = 8'h00;
    mem[490] = 8'h00;
    mem[491] = 8'h00;
    mem[492] = 8'h00;
    mem[493] = 8'h00;
    mem[494] = 8'h00;
    mem[495] = 8'h00;
    mem[496] = 8'h00;
    mem[497] = 8'h00;
    mem[498] = 8'h00;
    mem[499] = 8'h00;
    mem[500] = 8'h00;
    mem[501] = 8'h00;
    mem[502] = 8'h00;
    mem[503] = 8'h00;
    mem[504] = 8'h00;
    mem[505] = 8'h00;
    mem[506] = 8'h00;
    mem[507] = 8'h00;
    mem[508] = 8'h00;
    mem[509] = 8'h00;
    mem[510] = 8'h00;
    mem[511] = 8'h00;
  end

  wire [8:0] addr = {y[5:0], x[5:3]};
  assign pixel = mem[addr][x&7];

endmodule
