module byte_receiver_formal ();
endmodule
