module fsm_260_states(
    input clk,
    input rst_n,
    output reg [8:0] state
);

// State definitions
parameter s1   = 9'd0;
parameter s2   = 9'd1;
parameter s3   = 9'd2;
parameter s4   = 9'd3;
parameter s5   = 9'd4;
parameter s6   = 9'd5;
parameter s7   = 9'd6;
parameter s8   = 9'd7;
parameter s9   = 9'd8;
parameter s10  = 9'd9;
parameter s11  = 9'd10;
parameter s12  = 9'd11;
parameter s13  = 9'd12;
parameter s14  = 9'd13;
parameter s15  = 9'd14;
parameter s16  = 9'd15;
parameter s17  = 9'd16;
parameter s18  = 9'd17;
parameter s19  = 9'd18;
parameter s20  = 9'd19;
parameter s21  = 9'd20;
parameter s22  = 9'd21;
parameter s23  = 9'd22;
parameter s24  = 9'd23;
parameter s25  = 9'd24;
parameter s26  = 9'd25;
parameter s27  = 9'd26;
parameter s28  = 9'd27;
parameter s29  = 9'd28;
parameter s30  = 9'd29;
parameter s31  = 9'd30;
parameter s32  = 9'd31;
parameter s33  = 9'd32;
parameter s34  = 9'd33;
parameter s35  = 9'd34;
parameter s36  = 9'd35;
parameter s37  = 9'd36;
parameter s38  = 9'd37;
parameter s39  = 9'd38;
parameter s40  = 9'd39;
parameter s41  = 9'd40;
parameter s42  = 9'd41;
parameter s43  = 9'd42;
parameter s44  = 9'd43;
parameter s45  = 9'd44;
parameter s46  = 9'd45;
parameter s47  = 9'd46;
parameter s48  = 9'd47;
parameter s49  = 9'd48;
parameter s50  = 9'd49;
parameter s51  = 9'd50;
parameter s52  = 9'd51;
parameter s53  = 9'd52;
parameter s54  = 9'd53;
parameter s55  = 9'd54;
parameter s56  = 9'd55;
parameter s57  = 9'd56;
parameter s58  = 9'd57;
parameter s59  = 9'd58;
parameter s60  = 9'd59;
parameter s61  = 9'd60;
parameter s62  = 9'd61;
parameter s63  = 9'd62;
parameter s64  = 9'd63;
parameter s65  = 9'd64;
parameter s66  = 9'd65;
parameter s67  = 9'd66;
parameter s68  = 9'd67;
parameter s69  = 9'd68;
parameter s70  = 9'd69;
parameter s71  = 9'd70;
parameter s72  = 9'd71;
parameter s73  = 9'd72;
parameter s74  = 9'd73;
parameter s75  = 9'd74;
parameter s76  = 9'd75;
parameter s77  = 9'd76;
parameter s78  = 9'd77;
parameter s79  = 9'd78;
parameter s80  = 9'd79;
parameter s81  = 9'd80;
parameter s82  = 9'd81;
parameter s83  = 9'd82;
parameter s84  = 9'd83;
parameter s85  = 9'd84;
parameter s86  = 9'd85;
parameter s87  = 9'd86;
parameter s88  = 9'd87;
parameter s89  = 9'd88;
parameter s90  = 9'd89;
parameter s91  = 9'd90;
parameter s92  = 9'd91;
parameter s93  = 9'd92;
parameter s94  = 9'd93;
parameter s95  = 9'd94;
parameter s96  = 9'd95;
parameter s97  = 9'd96;
parameter s98  = 9'd97;
parameter s99  = 9'd98;
parameter s100 = 9'd99;
parameter s101 = 9'd100;
parameter s102 = 9'd101;
parameter s103 = 9'd102;
parameter s104 = 9'd103;
parameter s105 = 9'd104;
parameter s106 = 9'd105;
parameter s107 = 9'd106;
parameter s108 = 9'd107;
parameter s109 = 9'd108;
parameter s110 = 9'd109;
parameter s111 = 9'd110;
parameter s112 = 9'd111;
parameter s113 = 9'd112;
parameter s114 = 9'd113;
parameter s115 = 9'd114;
parameter s116 = 9'd115;
parameter s117 = 9'd116;
parameter s118 = 9'd117;
parameter s119 = 9'd118;
parameter s120 = 9'd119;
parameter s121 = 9'd120;
parameter s122 = 9'd121;
parameter s123 = 9'd122;
parameter s124 = 9'd123;
parameter s125 = 9'd124;
parameter s126 = 9'd125;
parameter s127 = 9'd126;
parameter s128 = 9'd127;
parameter s129 = 9'd128;
parameter s130 = 9'd129;
parameter s131 = 9'd130;
parameter s132 = 9'd131;
parameter s133 = 9'd132;
parameter s134 = 9'd133;
parameter s135 = 9'd134;
parameter s136 = 9'd135;
parameter s137 = 9'd136;
parameter s138 = 9'd137;
parameter s139 = 9'd138;
parameter s140 = 9'd139;
parameter s141 = 9'd140;
parameter s142 = 9'd141;
parameter s143 = 9'd142;
parameter s144 = 9'd143;
parameter s145 = 9'd144;
parameter s146 = 9'd145;
parameter s147 = 9'd146;
parameter s148 = 9'd147;
parameter s149 = 9'd148;
parameter s150 = 9'd149;
parameter s151 = 9'd150;
parameter s152 = 9'd151;
parameter s153 = 9'd152;
parameter s154 = 9'd153;
parameter s155 = 9'd154;
parameter s156 = 9'd155;
parameter s157 = 9'd156;
parameter s158 = 9'd157;
parameter s159 = 9'd158;
parameter s160 = 9'd159;
parameter s161 = 9'd160;
parameter s162 = 9'd161;
parameter s163 = 9'd162;
parameter s164 = 9'd163;
parameter s165 = 9'd164;
parameter s166 = 9'd165;
parameter s167 = 9'd166;
parameter s168 = 9'd167;
parameter s169 = 9'd168;
parameter s170 = 9'd169;
parameter s171 = 9'd170;
parameter s172 = 9'd171;
parameter s173 = 9'd172;
parameter s174 = 9'd173;
parameter s175 = 9'd174;
parameter s176 = 9'd175;
parameter s177 = 9'd176;
parameter s178 = 9'd177;
parameter s179 = 9'd178;
parameter s180 = 9'd179;
parameter s181 = 9'd180;
parameter s182 = 9'd181;
parameter s183 = 9'd182;
parameter s184 = 9'd183;
parameter s185 = 9'd184;
parameter s186 = 9'd185;
parameter s187 = 9'd186;
parameter s188 = 9'd187;
parameter s189 = 9'd188;
parameter s190 = 9'd189;
parameter s191 = 9'd190;
parameter s192 = 9'd191;
parameter s193 = 9'd192;
parameter s194 = 9'd193;
parameter s195 = 9'd194;
parameter s196 = 9'd195;
parameter s197 = 9'd196;
parameter s198 = 9'd197;
parameter s199 = 9'd198;
parameter s200 = 9'd199;
parameter s201 = 9'd200;
parameter s202 = 9'd201;
parameter s203 = 9'd202;
parameter s204 = 9'd203;
parameter s205 = 9'd204;
parameter s206 = 9'd205;
parameter s207 = 9'd206;
parameter s208 = 9'd207;
parameter s209 = 9'd208;
parameter s210 = 9'd209;
parameter s211 = 9'd210;
parameter s212 = 9'd211;
parameter s213 = 9'd212;
parameter s214 = 9'd213;
parameter s215 = 9'd214;
parameter s216 = 9'd215;
parameter s217 = 9'd216;
parameter s218 = 9'd217;
parameter s219 = 9'd218;
parameter s220 = 9'd219;
parameter s221 = 9'd220;
parameter s222 = 9'd221;
parameter s223 = 9'd222;
parameter s224 = 9'd223;
parameter s225 = 9'd224;
parameter s226 = 9'd225;
parameter s227 = 9'd226;
parameter s228 = 9'd227;
parameter s229 = 9'd228;
parameter s230 = 9'd229;
parameter s231 = 9'd230;
parameter s232 = 9'd231;
parameter s233 = 9'd232;
parameter s234 = 9'd233;
parameter s235 = 9'd234;
parameter s236 = 9'd235;
parameter s237 = 9'd236;
parameter s238 = 9'd237;
parameter s239 = 9'd238;
parameter s240 = 9'd239;
parameter s241 = 9'd240;
parameter s242 = 9'd241;
parameter s243 = 9'd242;
parameter s244 = 9'd243;
parameter s245 = 9'd244;
parameter s246 = 9'd245;
parameter s247 = 9'd246;
parameter s248 = 9'd247;
parameter s249 = 9'd248;
parameter s250 = 9'd249;
parameter s251 = 9'd250;
parameter s252 = 9'd251;
parameter s253 = 9'd252;
parameter s254 = 9'd253;
parameter s255 = 9'd254;
parameter s256 = 9'd255;
parameter s257 = 9'd256;
parameter s258 = 9'd257;
parameter s259 = 9'd258;
parameter s260 = 9'd259;



always @(posedge clk or negedge rst_n) begin
    if (!rst_n) begin
        state <= s1;
    end else begin
        case (state)
            s1: state <= s2;
            s2: state <= s3;
            s3: state <= s4;
            s4: state <= s5;
            s5: state <= s6;
            s6: state <= s7;
            s7: state <= s8;
            s8: state <= s9;
            s9: state <= s10;
            s10: state <= s11;
            s11: state <= s12;
            s12: state <= s13;
            s13: state <= s14;
            s14: state <= s15;
            s15: state <= s16;
            s16: state <= s17;
            s17: state <= s18;
            s18: state <= s19;
            s19: state <= s20;
            s20: state <= s21;
            s21: state <= s22;
            s22: state <= s23;
            s23: state <= s24;
            s24: state <= s25;
            s25: state <= s26;
            s26: state <= s27;
            s27: state <= s28;
            s28: state <= s29;
            s29: state <= s30;
            s30: state <= s31;
            s31: state <= s32;
            s32: state <= s33;
            s33: state <= s34;
            s34: state <= s35;
            s35: state <= s36;
            s36: state <= s37;
            s37: state <= s38;
            s38: state <= s39;
            s39: state <= s40;
            s40: state <= s41;
            s41: state <= s42;
            s42: state <= s43;
            s43: state <= s44;
            s44: state <= s45;
            s45: state <= s46;
            s46: state <= s47;
            s47: state <= s48;
            s48: state <= s49;
            s49: state <= s50;
            s50: state <= s51;
            s51: state <= s52;
            s52: state <= s53;
            s53: state <= s54;
            s54: state <= s55;
            s55: state <= s56;
            s56: state <= s57;
            s57: state <= s58;
            s58: state <= s59;
            s59: state <= s60;
            s60: state <= s61;
            s61: state <= s62;
            s62: state <= s63;
            s63: state <= s64;
            s64: state <= s65;
            s65: state <= s66;
            s66: state <= s67;
            s67: state <= s68;
            s68: state <= s69;
            s69: state <= s70;
            s70: state <= s71;
            s71: state <= s72;
            s72: state <= s73;
            s73: state <= s74;
            s74: state <= s75;
            s75: state <= s76;
            s76: state <= s77;
            s77: state <= s78;
            s78: state <= s79;
            s79: state <= s80;
            s80: state <= s81;
            s81: state <= s82;
            s82: state <= s83;
            s83: state <= s84;
            s84: state <= s85;
            s85: state <= s86;
            s86: state <= s87;
            s87: state <= s88;
            s88: state <= s89;
            s89: state <= s90;
            s90: state <= s91;
            s91: state <= s92;
            s92: state <= s93;
            s93: state <= s94;
            s94: state <= s95;
            s95: state <= s96;
            s96: state <= s97;
            s97: state <= s98;
            s98: state <= s99;
            s99: state <= s100;
            s100: state <= s101;
            s101: state <= s102;
            s102: state <= s103;
            s103: state <= s104;
            s104: state <= s105;
            s105: state <= s106;
            s106: state <= s107;
            s107: state <= s108;
            s108: state <= s109;
            s109: state <= s110;
            s110: state <= s111;
            s111: state <= s112;
            s112: state <= s113;
            s113: state <= s114;
            s114: state <= s115;
            s115: state <= s116;
            s116: state <= s117;
            s117: state <= s118;
            s118: state <= s119;
            s119: state <= s120;
            s120: state <= s121;
            s121: state <= s122;
            s122: state <= s123;
            s123: state <= s124;
            s124: state <= s125;
            s125: state <= s126;
            s126: state <= s127;
            s127: state <= s128;
            s128: state <= s129;
            s129: state <= s130;
            s130: state <= s131;
            s131: state <= s132;
            s132: state <= s133;
            s133: state <= s134;
            s134: state <= s135;
            s135: state <= s136;
            s136: state <= s137;
            s137: state <= s138;
            s138: state <= s139;
            s139: state <= s140;
            s140: state <= s141;
            s141: state <= s142;
            s142: state <= s143;
            s143: state <= s144;
            s144: state <= s145;
            s145: state <= s146;
            s146: state <= s147;
            s147: state <= s148;
            s148: state <= s149;
            s149: state <= s150;
            s150: state <= s151;
            s151: state <= s152;
            s152: state <= s153;
            s153: state <= s154;
            s154: state <= s155;
            s155: state <= s156;
            s156: state <= s157;
            s157: state <= s158;
            s158: state <= s159;
            s159: state <= s160;
            s160: state <= s161;
            s161: state <= s162;
            s162: state <= s163;
            s163: state <= s164;
            s164: state <= s165;
            s165: state <= s166;
            s166: state <= s167;
            s167: state <= s168;
            s168: state <= s169;
            s169: state <= s170;
            s170: state <= s171;
            s171: state <= s172;
            s172: state <= s173;
            s173: state <= s174;
            s174: state <= s175;
            s175: state <= s176;
            s176: state <= s177;
            s177: state <= s178;
            s178: state <= s179;
            s179: state <= s180;
            s180: state <= s181;
            s181: state <= s182;
            s182: state <= s183;
            s183: state <= s184;
            s184: state <= s185;
            s185: state <= s186;
            s186: state <= s187;
            s187: state <= s188;
            s188: state <= s189;
            s189: state <= s190;
            s190: state <= s191;
            s191: state <= s192;
            s192: state <= s193;
            s193: state <= s194;
            s194: state <= s195;
            s195: state <= s196;
            s196: state <= s197;
            s197: state <= s198;
            s198: state <= s199;
            s199: state <= s200;
            s200: state <= s201;
            s201: state <= s202;
            s202: state <= s203;
            s203: state <= s204;
            s204: state <= s205;
            s205: state <= s206;
            s206: state <= s207;
            s207: state <= s208;
            s208: state <= s209;
            s209: state <= s210;
            s210: state <= s211;
            s211: state <= s212;
            s212: state <= s213;
            s213: state <= s214;
            s214: state <= s215;
            s215: state <= s216;
            s216: state <= s217;
            s217: state <= s218;
            s218: state <= s219;
            s219: state <= s220;
            s220: state <= s221;
            s221: state <= s222;
            s222: state <= s223;
            s223: state <= s224;
            s224: state <= s225;
            s225: state <= s226;
            s226: state <= s227;
            s227: state <= s228;
            s228: state <= s229;
            s229: state <= s230;
            s230: state <= s231;
            s231: state <= s232;
            s232: state <= s233;
            s233: state <= s234;
            s234: state <= s235;
            s235: state <= s236;
            s236: state <= s237;
            s237: state <= s238;
            s238: state <= s239;
            s239: state <= s240;
            s240: state <= s241;
            s241: state <= s242;
            s242: state <= s243;
            s243: state <= s244;
            s244: state <= s245;
            s245: state <= s246;
            s246: state <= s247;
            s247: state <= s248;
            s248: state <= s249;
            s249: state <= s250;
            s250: state <= s251;
            s251: state <= s252;
            s252: state <= s253;
            s253: state <= s254;
            s254: state <= s255;
            s255: state <= s256;
            s256: state <= s257;
            s257: state <= s258;
            s258: state <= s259;
            //s259: state <= s1;
            s259: state <= s260;
            s260: state <= s1; // or another state as needed

            default: begin
                // Handle any unexpected states
                state <= s1; // or some error state
            end
        endcase
    end
end

endmodule
