module logo_table(
		input wire [11:0] addr,
		output wire data
	);

	reg d;
	always @(*) begin
		case (addr)
			0: d = 0;
			1: d = 0;
			2: d = 0;
			3: d = 0;
			4: d = 0;
			5: d = 0;
			6: d = 0;
			7: d = 0;
			8: d = 1;
			9: d = 0;
			10: d = 1;
			11: d = 1;
			12: d = 1;
			13: d = 1;
			14: d = 0;
			15: d = 0;
			16: d = 0;
			17: d = 0;
			18: d = 0;
			19: d = 0;
			20: d = 0;
			21: d = 0;
			22: d = 0;
			23: d = 0;
			24: d = 0;
			25: d = 0;
			26: d = 0;
			27: d = 0;
			28: d = 1;
			29: d = 0;
			30: d = 0;
			31: d = 0;
			32: d = 0;
			33: d = 0;
			34: d = 0;
			35: d = 0;
			36: d = 0;
			37: d = 0;
			38: d = 0;
			39: d = 0;
			40: d = 0;
			41: d = 0;
			42: d = 0;
			43: d = 0;
			44: d = 0;
			45: d = 0;
			46: d = 0;
			47: d = 0;
			48: d = 0;
			49: d = 0;
			50: d = 0;
			51: d = 0;
			52: d = 0;
			53: d = 0;
			54: d = 0;
			55: d = 0;
			56: d = 0;
			57: d = 0;
			58: d = 0;
			59: d = 0;
			60: d = 0;
			61: d = 0;
			62: d = 0;
			63: d = 0;
			64: d = 0;
			65: d = 0;
			66: d = 0;
			67: d = 0;
			68: d = 0;
			69: d = 0;
			70: d = 0;
			71: d = 0;
			72: d = 0;
			73: d = 0;
			74: d = 0;
			75: d = 0;
			76: d = 0;
			77: d = 0;
			78: d = 0;
			79: d = 0;
			80: d = 0;
			81: d = 0;
			82: d = 0;
			83: d = 0;
			84: d = 0;
			85: d = 0;
			86: d = 0;
			87: d = 0;
			88: d = 0;
			89: d = 0;
			90: d = 0;
			91: d = 0;
			92: d = 0;
			93: d = 0;
			94: d = 0;
			95: d = 0;
			96: d = 0;
			97: d = 0;
			98: d = 0;
			99: d = 0;
			100: d = 0;
			101: d = 0;
			102: d = 0;
			103: d = 0;
			104: d = 0;
			105: d = 0;
			106: d = 0;
			107: d = 0;
			108: d = 0;
			109: d = 0;
			110: d = 0;
			111: d = 0;
			112: d = 0;
			113: d = 0;
			114: d = 0;
			115: d = 0;
			116: d = 0;
			117: d = 0;
			118: d = 0;
			119: d = 0;
			120: d = 0;
			121: d = 0;
			122: d = 0;
			123: d = 0;
			124: d = 0;
			125: d = 0;
			126: d = 0;
			127: d = 0;
			128: d = 0;
			129: d = 0;
			130: d = 0;
			131: d = 0;
			132: d = 0;
			133: d = 0;
			134: d = 1;
			135: d = 0;
			136: d = 0;
			137: d = 0;
			138: d = 1;
			139: d = 0;
			140: d = 0;
			141: d = 1;
			142: d = 0;
			143: d = 0;
			144: d = 0;
			145: d = 0;
			146: d = 0;
			147: d = 0;
			148: d = 0;
			149: d = 0;
			150: d = 0;
			151: d = 0;
			152: d = 0;
			153: d = 0;
			154: d = 1;
			155: d = 0;
			156: d = 1;
			157: d = 1;
			158: d = 0;
			159: d = 0;
			160: d = 0;
			161: d = 0;
			162: d = 0;
			163: d = 0;
			164: d = 0;
			165: d = 0;
			166: d = 0;
			167: d = 0;
			168: d = 0;
			169: d = 0;
			170: d = 0;
			171: d = 0;
			172: d = 0;
			173: d = 0;
			174: d = 0;
			175: d = 0;
			176: d = 0;
			177: d = 0;
			178: d = 0;
			179: d = 0;
			180: d = 0;
			181: d = 0;
			182: d = 0;
			183: d = 0;
			184: d = 0;
			185: d = 0;
			186: d = 0;
			187: d = 0;
			188: d = 0;
			189: d = 0;
			190: d = 0;
			191: d = 0;
			192: d = 0;
			193: d = 0;
			194: d = 0;
			195: d = 0;
			196: d = 0;
			197: d = 0;
			198: d = 0;
			199: d = 0;
			200: d = 0;
			201: d = 0;
			202: d = 0;
			203: d = 0;
			204: d = 0;
			205: d = 0;
			206: d = 0;
			207: d = 0;
			208: d = 0;
			209: d = 0;
			210: d = 0;
			211: d = 0;
			212: d = 0;
			213: d = 0;
			214: d = 0;
			215: d = 0;
			216: d = 0;
			217: d = 0;
			218: d = 0;
			219: d = 0;
			220: d = 0;
			221: d = 0;
			222: d = 0;
			223: d = 0;
			224: d = 0;
			225: d = 0;
			226: d = 0;
			227: d = 0;
			228: d = 0;
			229: d = 0;
			230: d = 0;
			231: d = 0;
			232: d = 0;
			233: d = 0;
			234: d = 0;
			235: d = 0;
			236: d = 0;
			237: d = 0;
			238: d = 0;
			239: d = 0;
			240: d = 0;
			241: d = 0;
			242: d = 0;
			243: d = 0;
			244: d = 0;
			245: d = 0;
			246: d = 0;
			247: d = 0;
			248: d = 0;
			249: d = 0;
			250: d = 0;
			251: d = 0;
			252: d = 0;
			253: d = 0;
			254: d = 0;
			255: d = 0;
			256: d = 0;
			257: d = 0;
			258: d = 0;
			259: d = 0;
			260: d = 1;
			261: d = 0;
			262: d = 1;
			263: d = 1;
			264: d = 1;
			265: d = 0;
			266: d = 0;
			267: d = 1;
			268: d = 1;
			269: d = 0;
			270: d = 0;
			271: d = 0;
			272: d = 0;
			273: d = 0;
			274: d = 0;
			275: d = 0;
			276: d = 0;
			277: d = 0;
			278: d = 0;
			279: d = 0;
			280: d = 1;
			281: d = 0;
			282: d = 1;
			283: d = 1;
			284: d = 1;
			285: d = 1;
			286: d = 0;
			287: d = 0;
			288: d = 0;
			289: d = 0;
			290: d = 0;
			291: d = 0;
			292: d = 0;
			293: d = 0;
			294: d = 0;
			295: d = 0;
			296: d = 0;
			297: d = 0;
			298: d = 0;
			299: d = 0;
			300: d = 0;
			301: d = 0;
			302: d = 0;
			303: d = 0;
			304: d = 0;
			305: d = 0;
			306: d = 0;
			307: d = 0;
			308: d = 0;
			309: d = 0;
			310: d = 0;
			311: d = 0;
			312: d = 0;
			313: d = 0;
			314: d = 0;
			315: d = 0;
			316: d = 0;
			317: d = 0;
			318: d = 0;
			319: d = 0;
			320: d = 0;
			321: d = 0;
			322: d = 0;
			323: d = 0;
			324: d = 0;
			325: d = 0;
			326: d = 0;
			327: d = 0;
			328: d = 0;
			329: d = 0;
			330: d = 0;
			331: d = 0;
			332: d = 0;
			333: d = 0;
			334: d = 0;
			335: d = 0;
			336: d = 0;
			337: d = 0;
			338: d = 0;
			339: d = 0;
			340: d = 0;
			341: d = 0;
			342: d = 0;
			343: d = 0;
			344: d = 0;
			345: d = 0;
			346: d = 0;
			347: d = 0;
			348: d = 0;
			349: d = 0;
			350: d = 0;
			351: d = 0;
			352: d = 0;
			353: d = 0;
			354: d = 0;
			355: d = 0;
			356: d = 0;
			357: d = 0;
			358: d = 0;
			359: d = 0;
			360: d = 0;
			361: d = 0;
			362: d = 0;
			363: d = 0;
			364: d = 1;
			365: d = 0;
			366: d = 1;
			367: d = 1;
			368: d = 0;
			369: d = 0;
			370: d = 0;
			371: d = 0;
			372: d = 0;
			373: d = 0;
			374: d = 0;
			375: d = 0;
			376: d = 0;
			377: d = 0;
			378: d = 0;
			379: d = 0;
			380: d = 0;
			381: d = 0;
			382: d = 0;
			383: d = 0;
			384: d = 0;
			385: d = 0;
			386: d = 1;
			387: d = 0;
			388: d = 0;
			389: d = 1;
			390: d = 1;
			391: d = 1;
			392: d = 0;
			393: d = 1;
			394: d = 1;
			395: d = 0;
			396: d = 1;
			397: d = 1;
			398: d = 0;
			399: d = 0;
			400: d = 0;
			401: d = 0;
			402: d = 0;
			403: d = 0;
			404: d = 0;
			405: d = 0;
			406: d = 1;
			407: d = 0;
			408: d = 0;
			409: d = 0;
			410: d = 1;
			411: d = 0;
			412: d = 0;
			413: d = 1;
			414: d = 0;
			415: d = 0;
			416: d = 0;
			417: d = 0;
			418: d = 0;
			419: d = 0;
			420: d = 0;
			421: d = 0;
			422: d = 0;
			423: d = 0;
			424: d = 0;
			425: d = 0;
			426: d = 0;
			427: d = 0;
			428: d = 0;
			429: d = 0;
			430: d = 0;
			431: d = 0;
			432: d = 0;
			433: d = 0;
			434: d = 0;
			435: d = 0;
			436: d = 0;
			437: d = 0;
			438: d = 0;
			439: d = 0;
			440: d = 0;
			441: d = 0;
			442: d = 0;
			443: d = 0;
			444: d = 0;
			445: d = 0;
			446: d = 0;
			447: d = 0;
			448: d = 0;
			449: d = 0;
			450: d = 0;
			451: d = 0;
			452: d = 0;
			453: d = 0;
			454: d = 0;
			455: d = 0;
			456: d = 0;
			457: d = 0;
			458: d = 0;
			459: d = 0;
			460: d = 0;
			461: d = 0;
			462: d = 0;
			463: d = 0;
			464: d = 0;
			465: d = 0;
			466: d = 0;
			467: d = 0;
			468: d = 0;
			469: d = 0;
			470: d = 0;
			471: d = 0;
			472: d = 0;
			473: d = 0;
			474: d = 0;
			475: d = 0;
			476: d = 0;
			477: d = 0;
			478: d = 0;
			479: d = 0;
			480: d = 0;
			481: d = 0;
			482: d = 0;
			483: d = 0;
			484: d = 0;
			485: d = 0;
			486: d = 0;
			487: d = 0;
			488: d = 0;
			489: d = 0;
			490: d = 1;
			491: d = 0;
			492: d = 0;
			493: d = 1;
			494: d = 0;
			495: d = 0;
			496: d = 0;
			497: d = 0;
			498: d = 0;
			499: d = 0;
			500: d = 0;
			501: d = 0;
			502: d = 0;
			503: d = 0;
			504: d = 0;
			505: d = 0;
			506: d = 0;
			507: d = 0;
			508: d = 0;
			509: d = 0;
			510: d = 0;
			511: d = 0;
			512: d = 0;
			513: d = 0;
			514: d = 1;
			515: d = 1;
			516: d = 0;
			517: d = 0;
			518: d = 0;
			519: d = 0;
			520: d = 1;
			521: d = 0;
			522: d = 0;
			523: d = 1;
			524: d = 0;
			525: d = 1;
			526: d = 0;
			527: d = 0;
			528: d = 0;
			529: d = 0;
			530: d = 0;
			531: d = 0;
			532: d = 1;
			533: d = 0;
			534: d = 1;
			535: d = 1;
			536: d = 1;
			537: d = 0;
			538: d = 0;
			539: d = 1;
			540: d = 1;
			541: d = 0;
			542: d = 0;
			543: d = 0;
			544: d = 0;
			545: d = 0;
			546: d = 0;
			547: d = 0;
			548: d = 0;
			549: d = 0;
			550: d = 0;
			551: d = 0;
			552: d = 0;
			553: d = 0;
			554: d = 0;
			555: d = 0;
			556: d = 0;
			557: d = 0;
			558: d = 0;
			559: d = 0;
			560: d = 0;
			561: d = 0;
			562: d = 0;
			563: d = 0;
			564: d = 0;
			565: d = 0;
			566: d = 0;
			567: d = 0;
			568: d = 0;
			569: d = 0;
			570: d = 0;
			571: d = 0;
			572: d = 0;
			573: d = 0;
			574: d = 0;
			575: d = 0;
			576: d = 0;
			577: d = 0;
			578: d = 0;
			579: d = 0;
			580: d = 0;
			581: d = 0;
			582: d = 0;
			583: d = 0;
			584: d = 0;
			585: d = 0;
			586: d = 0;
			587: d = 0;
			588: d = 0;
			589: d = 0;
			590: d = 0;
			591: d = 0;
			592: d = 0;
			593: d = 0;
			594: d = 0;
			595: d = 0;
			596: d = 0;
			597: d = 0;
			598: d = 0;
			599: d = 0;
			600: d = 0;
			601: d = 0;
			602: d = 0;
			603: d = 0;
			604: d = 0;
			605: d = 0;
			606: d = 0;
			607: d = 0;
			608: d = 0;
			609: d = 0;
			610: d = 0;
			611: d = 0;
			612: d = 0;
			613: d = 0;
			614: d = 0;
			615: d = 0;
			616: d = 0;
			617: d = 0;
			618: d = 1;
			619: d = 1;
			620: d = 1;
			621: d = 0;
			622: d = 0;
			623: d = 1;
			624: d = 0;
			625: d = 0;
			626: d = 0;
			627: d = 0;
			628: d = 0;
			629: d = 0;
			630: d = 0;
			631: d = 0;
			632: d = 0;
			633: d = 0;
			634: d = 0;
			635: d = 0;
			636: d = 0;
			637: d = 0;
			638: d = 0;
			639: d = 0;
			640: d = 0;
			641: d = 0;
			642: d = 1;
			643: d = 1;
			644: d = 0;
			645: d = 1;
			646: d = 1;
			647: d = 0;
			648: d = 1;
			649: d = 1;
			650: d = 0;
			651: d = 0;
			652: d = 0;
			653: d = 0;
			654: d = 0;
			655: d = 0;
			656: d = 0;
			657: d = 0;
			658: d = 1;
			659: d = 0;
			660: d = 0;
			661: d = 1;
			662: d = 1;
			663: d = 1;
			664: d = 0;
			665: d = 1;
			666: d = 1;
			667: d = 0;
			668: d = 0;
			669: d = 1;
			670: d = 0;
			671: d = 0;
			672: d = 0;
			673: d = 0;
			674: d = 0;
			675: d = 0;
			676: d = 0;
			677: d = 0;
			678: d = 0;
			679: d = 0;
			680: d = 0;
			681: d = 0;
			682: d = 0;
			683: d = 0;
			684: d = 0;
			685: d = 0;
			686: d = 0;
			687: d = 0;
			688: d = 0;
			689: d = 0;
			690: d = 0;
			691: d = 0;
			692: d = 0;
			693: d = 0;
			694: d = 0;
			695: d = 0;
			696: d = 0;
			697: d = 0;
			698: d = 0;
			699: d = 0;
			700: d = 0;
			701: d = 0;
			702: d = 0;
			703: d = 0;
			704: d = 0;
			705: d = 0;
			706: d = 0;
			707: d = 0;
			708: d = 0;
			709: d = 0;
			710: d = 0;
			711: d = 0;
			712: d = 0;
			713: d = 0;
			714: d = 0;
			715: d = 0;
			716: d = 0;
			717: d = 0;
			718: d = 0;
			719: d = 0;
			720: d = 0;
			721: d = 0;
			722: d = 0;
			723: d = 0;
			724: d = 0;
			725: d = 0;
			726: d = 0;
			727: d = 0;
			728: d = 0;
			729: d = 0;
			730: d = 0;
			731: d = 0;
			732: d = 0;
			733: d = 0;
			734: d = 0;
			735: d = 0;
			736: d = 0;
			737: d = 0;
			738: d = 0;
			739: d = 0;
			740: d = 0;
			741: d = 0;
			742: d = 0;
			743: d = 0;
			744: d = 0;
			745: d = 0;
			746: d = 1;
			747: d = 1;
			748: d = 0;
			749: d = 1;
			750: d = 0;
			751: d = 0;
			752: d = 0;
			753: d = 0;
			754: d = 0;
			755: d = 0;
			756: d = 0;
			757: d = 0;
			758: d = 0;
			759: d = 0;
			760: d = 0;
			761: d = 0;
			762: d = 0;
			763: d = 0;
			764: d = 0;
			765: d = 0;
			766: d = 0;
			767: d = 0;
			768: d = 0;
			769: d = 0;
			770: d = 0;
			771: d = 1;
			772: d = 1;
			773: d = 0;
			774: d = 0;
			775: d = 1;
			776: d = 0;
			777: d = 1;
			778: d = 1;
			779: d = 0;
			780: d = 1;
			781: d = 1;
			782: d = 0;
			783: d = 0;
			784: d = 0;
			785: d = 0;
			786: d = 1;
			787: d = 1;
			788: d = 0;
			789: d = 0;
			790: d = 0;
			791: d = 0;
			792: d = 1;
			793: d = 0;
			794: d = 0;
			795: d = 1;
			796: d = 1;
			797: d = 0;
			798: d = 0;
			799: d = 0;
			800: d = 0;
			801: d = 0;
			802: d = 0;
			803: d = 0;
			804: d = 0;
			805: d = 0;
			806: d = 0;
			807: d = 0;
			808: d = 0;
			809: d = 0;
			810: d = 1;
			811: d = 0;
			812: d = 1;
			813: d = 1;
			814: d = 0;
			815: d = 0;
			816: d = 0;
			817: d = 0;
			818: d = 0;
			819: d = 0;
			820: d = 0;
			821: d = 0;
			822: d = 0;
			823: d = 0;
			824: d = 0;
			825: d = 0;
			826: d = 0;
			827: d = 0;
			828: d = 0;
			829: d = 0;
			830: d = 0;
			831: d = 0;
			832: d = 0;
			833: d = 0;
			834: d = 0;
			835: d = 0;
			836: d = 0;
			837: d = 0;
			838: d = 0;
			839: d = 0;
			840: d = 0;
			841: d = 0;
			842: d = 0;
			843: d = 0;
			844: d = 0;
			845: d = 0;
			846: d = 0;
			847: d = 0;
			848: d = 0;
			849: d = 0;
			850: d = 0;
			851: d = 0;
			852: d = 0;
			853: d = 0;
			854: d = 0;
			855: d = 0;
			856: d = 0;
			857: d = 0;
			858: d = 0;
			859: d = 0;
			860: d = 0;
			861: d = 0;
			862: d = 0;
			863: d = 0;
			864: d = 0;
			865: d = 0;
			866: d = 0;
			867: d = 0;
			868: d = 0;
			869: d = 0;
			870: d = 0;
			871: d = 0;
			872: d = 0;
			873: d = 0;
			874: d = 1;
			875: d = 1;
			876: d = 1;
			877: d = 0;
			878: d = 0;
			879: d = 1;
			880: d = 0;
			881: d = 0;
			882: d = 0;
			883: d = 0;
			884: d = 0;
			885: d = 0;
			886: d = 0;
			887: d = 0;
			888: d = 0;
			889: d = 0;
			890: d = 0;
			891: d = 0;
			892: d = 0;
			893: d = 0;
			894: d = 0;
			895: d = 0;
			896: d = 0;
			897: d = 0;
			898: d = 0;
			899: d = 0;
			900: d = 1;
			901: d = 1;
			902: d = 0;
			903: d = 0;
			904: d = 1;
			905: d = 0;
			906: d = 0;
			907: d = 1;
			908: d = 1;
			909: d = 1;
			910: d = 0;
			911: d = 0;
			912: d = 0;
			913: d = 0;
			914: d = 1;
			915: d = 1;
			916: d = 0;
			917: d = 1;
			918: d = 1;
			919: d = 0;
			920: d = 1;
			921: d = 1;
			922: d = 1;
			923: d = 0;
			924: d = 0;
			925: d = 1;
			926: d = 0;
			927: d = 0;
			928: d = 0;
			929: d = 0;
			930: d = 0;
			931: d = 0;
			932: d = 0;
			933: d = 0;
			934: d = 0;
			935: d = 0;
			936: d = 1;
			937: d = 0;
			938: d = 0;
			939: d = 1;
			940: d = 0;
			941: d = 1;
			942: d = 0;
			943: d = 0;
			944: d = 0;
			945: d = 0;
			946: d = 0;
			947: d = 0;
			948: d = 0;
			949: d = 0;
			950: d = 0;
			951: d = 0;
			952: d = 0;
			953: d = 0;
			954: d = 0;
			955: d = 0;
			956: d = 0;
			957: d = 0;
			958: d = 0;
			959: d = 0;
			960: d = 0;
			961: d = 0;
			962: d = 0;
			963: d = 0;
			964: d = 0;
			965: d = 0;
			966: d = 0;
			967: d = 0;
			968: d = 0;
			969: d = 0;
			970: d = 0;
			971: d = 0;
			972: d = 0;
			973: d = 0;
			974: d = 0;
			975: d = 0;
			976: d = 1;
			977: d = 0;
			978: d = 0;
			979: d = 0;
			980: d = 0;
			981: d = 0;
			982: d = 0;
			983: d = 0;
			984: d = 0;
			985: d = 0;
			986: d = 0;
			987: d = 0;
			988: d = 0;
			989: d = 0;
			990: d = 0;
			991: d = 0;
			992: d = 0;
			993: d = 0;
			994: d = 0;
			995: d = 0;
			996: d = 0;
			997: d = 0;
			998: d = 0;
			999: d = 0;
			1000: d = 0;
			1001: d = 0;
			1002: d = 1;
			1003: d = 1;
			1004: d = 0;
			1005: d = 1;
			1006: d = 0;
			1007: d = 0;
			1008: d = 0;
			1009: d = 0;
			1010: d = 0;
			1011: d = 0;
			1012: d = 0;
			1013: d = 0;
			1014: d = 0;
			1015: d = 0;
			1016: d = 0;
			1017: d = 0;
			1018: d = 0;
			1019: d = 0;
			1020: d = 0;
			1021: d = 0;
			1022: d = 0;
			1023: d = 0;
			1024: d = 0;
			1025: d = 0;
			1026: d = 0;
			1027: d = 0;
			1028: d = 0;
			1029: d = 1;
			1030: d = 1;
			1031: d = 0;
			1032: d = 0;
			1033: d = 1;
			1034: d = 1;
			1035: d = 1;
			1036: d = 1;
			1037: d = 1;
			1038: d = 0;
			1039: d = 0;
			1040: d = 0;
			1041: d = 0;
			1042: d = 0;
			1043: d = 1;
			1044: d = 1;
			1045: d = 0;
			1046: d = 0;
			1047: d = 1;
			1048: d = 1;
			1049: d = 1;
			1050: d = 0;
			1051: d = 1;
			1052: d = 1;
			1053: d = 0;
			1054: d = 0;
			1055: d = 0;
			1056: d = 0;
			1057: d = 0;
			1058: d = 0;
			1059: d = 0;
			1060: d = 0;
			1061: d = 0;
			1062: d = 0;
			1063: d = 0;
			1064: d = 1;
			1065: d = 1;
			1066: d = 0;
			1067: d = 0;
			1068: d = 0;
			1069: d = 0;
			1070: d = 0;
			1071: d = 0;
			1072: d = 0;
			1073: d = 0;
			1074: d = 0;
			1075: d = 0;
			1076: d = 0;
			1077: d = 0;
			1078: d = 0;
			1079: d = 0;
			1080: d = 0;
			1081: d = 0;
			1082: d = 0;
			1083: d = 0;
			1084: d = 0;
			1085: d = 0;
			1086: d = 0;
			1087: d = 0;
			1088: d = 0;
			1089: d = 0;
			1090: d = 0;
			1091: d = 0;
			1092: d = 0;
			1093: d = 0;
			1094: d = 0;
			1095: d = 0;
			1096: d = 0;
			1097: d = 0;
			1098: d = 0;
			1099: d = 0;
			1100: d = 0;
			1101: d = 0;
			1102: d = 0;
			1103: d = 0;
			1104: d = 1;
			1105: d = 1;
			1106: d = 0;
			1107: d = 0;
			1108: d = 0;
			1109: d = 0;
			1110: d = 0;
			1111: d = 0;
			1112: d = 0;
			1113: d = 0;
			1114: d = 0;
			1115: d = 0;
			1116: d = 0;
			1117: d = 0;
			1118: d = 0;
			1119: d = 0;
			1120: d = 0;
			1121: d = 0;
			1122: d = 0;
			1123: d = 0;
			1124: d = 0;
			1125: d = 0;
			1126: d = 0;
			1127: d = 0;
			1128: d = 0;
			1129: d = 0;
			1130: d = 0;
			1131: d = 0;
			1132: d = 1;
			1133: d = 0;
			1134: d = 1;
			1135: d = 1;
			1136: d = 0;
			1137: d = 0;
			1138: d = 0;
			1139: d = 0;
			1140: d = 0;
			1141: d = 0;
			1142: d = 0;
			1143: d = 0;
			1144: d = 0;
			1145: d = 0;
			1146: d = 0;
			1147: d = 0;
			1148: d = 0;
			1149: d = 0;
			1150: d = 0;
			1151: d = 0;
			1152: d = 0;
			1153: d = 0;
			1154: d = 0;
			1155: d = 0;
			1156: d = 1;
			1157: d = 0;
			1158: d = 0;
			1159: d = 1;
			1160: d = 1;
			1161: d = 0;
			1162: d = 0;
			1163: d = 1;
			1164: d = 0;
			1165: d = 0;
			1166: d = 0;
			1167: d = 0;
			1168: d = 0;
			1169: d = 0;
			1170: d = 0;
			1171: d = 0;
			1172: d = 0;
			1173: d = 1;
			1174: d = 1;
			1175: d = 0;
			1176: d = 0;
			1177: d = 1;
			1178: d = 1;
			1179: d = 0;
			1180: d = 0;
			1181: d = 1;
			1182: d = 0;
			1183: d = 0;
			1184: d = 0;
			1185: d = 0;
			1186: d = 0;
			1187: d = 0;
			1188: d = 0;
			1189: d = 0;
			1190: d = 0;
			1191: d = 0;
			1192: d = 0;
			1193: d = 1;
			1194: d = 1;
			1195: d = 0;
			1196: d = 1;
			1197: d = 1;
			1198: d = 0;
			1199: d = 0;
			1200: d = 0;
			1201: d = 0;
			1202: d = 0;
			1203: d = 0;
			1204: d = 0;
			1205: d = 0;
			1206: d = 0;
			1207: d = 0;
			1208: d = 1;
			1209: d = 0;
			1210: d = 1;
			1211: d = 1;
			1212: d = 0;
			1213: d = 0;
			1214: d = 0;
			1215: d = 0;
			1216: d = 0;
			1217: d = 0;
			1218: d = 0;
			1219: d = 0;
			1220: d = 0;
			1221: d = 0;
			1222: d = 0;
			1223: d = 0;
			1224: d = 0;
			1225: d = 0;
			1226: d = 0;
			1227: d = 0;
			1228: d = 0;
			1229: d = 0;
			1230: d = 0;
			1231: d = 0;
			1232: d = 1;
			1233: d = 1;
			1234: d = 0;
			1235: d = 0;
			1236: d = 0;
			1237: d = 0;
			1238: d = 0;
			1239: d = 0;
			1240: d = 1;
			1241: d = 0;
			1242: d = 1;
			1243: d = 1;
			1244: d = 0;
			1245: d = 0;
			1246: d = 0;
			1247: d = 0;
			1248: d = 0;
			1249: d = 0;
			1250: d = 0;
			1251: d = 0;
			1252: d = 0;
			1253: d = 0;
			1254: d = 0;
			1255: d = 0;
			1256: d = 0;
			1257: d = 0;
			1258: d = 1;
			1259: d = 0;
			1260: d = 0;
			1261: d = 1;
			1262: d = 1;
			1263: d = 1;
			1264: d = 0;
			1265: d = 0;
			1266: d = 0;
			1267: d = 0;
			1268: d = 0;
			1269: d = 0;
			1270: d = 0;
			1271: d = 0;
			1272: d = 1;
			1273: d = 0;
			1274: d = 1;
			1275: d = 1;
			1276: d = 0;
			1277: d = 0;
			1278: d = 0;
			1279: d = 0;
			1280: d = 0;
			1281: d = 0;
			1282: d = 0;
			1283: d = 0;
			1284: d = 1;
			1285: d = 1;
			1286: d = 1;
			1287: d = 1;
			1288: d = 0;
			1289: d = 1;
			1290: d = 1;
			1291: d = 0;
			1292: d = 1;
			1293: d = 1;
			1294: d = 0;
			1295: d = 0;
			1296: d = 0;
			1297: d = 0;
			1298: d = 0;
			1299: d = 0;
			1300: d = 1;
			1301: d = 0;
			1302: d = 0;
			1303: d = 1;
			1304: d = 1;
			1305: d = 0;
			1306: d = 1;
			1307: d = 1;
			1308: d = 1;
			1309: d = 1;
			1310: d = 0;
			1311: d = 0;
			1312: d = 0;
			1313: d = 0;
			1314: d = 0;
			1315: d = 0;
			1316: d = 0;
			1317: d = 0;
			1318: d = 0;
			1319: d = 0;
			1320: d = 1;
			1321: d = 0;
			1322: d = 0;
			1323: d = 1;
			1324: d = 1;
			1325: d = 1;
			1326: d = 0;
			1327: d = 0;
			1328: d = 0;
			1329: d = 0;
			1330: d = 0;
			1331: d = 0;
			1332: d = 0;
			1333: d = 0;
			1334: d = 1;
			1335: d = 0;
			1336: d = 0;
			1337: d = 1;
			1338: d = 0;
			1339: d = 1;
			1340: d = 0;
			1341: d = 0;
			1342: d = 0;
			1343: d = 0;
			1344: d = 0;
			1345: d = 0;
			1346: d = 0;
			1347: d = 0;
			1348: d = 0;
			1349: d = 0;
			1350: d = 0;
			1351: d = 0;
			1352: d = 0;
			1353: d = 0;
			1354: d = 1;
			1355: d = 0;
			1356: d = 1;
			1357: d = 1;
			1358: d = 1;
			1359: d = 0;
			1360: d = 0;
			1361: d = 1;
			1362: d = 0;
			1363: d = 0;
			1364: d = 0;
			1365: d = 0;
			1366: d = 1;
			1367: d = 0;
			1368: d = 0;
			1369: d = 1;
			1370: d = 0;
			1371: d = 1;
			1372: d = 0;
			1373: d = 0;
			1374: d = 0;
			1375: d = 0;
			1376: d = 0;
			1377: d = 0;
			1378: d = 0;
			1379: d = 0;
			1380: d = 0;
			1381: d = 0;
			1382: d = 0;
			1383: d = 0;
			1384: d = 0;
			1385: d = 0;
			1386: d = 0;
			1387: d = 1;
			1388: d = 1;
			1389: d = 0;
			1390: d = 0;
			1391: d = 1;
			1392: d = 0;
			1393: d = 0;
			1394: d = 0;
			1395: d = 0;
			1396: d = 0;
			1397: d = 0;
			1398: d = 1;
			1399: d = 0;
			1400: d = 0;
			1401: d = 1;
			1402: d = 0;
			1403: d = 1;
			1404: d = 0;
			1405: d = 0;
			1406: d = 0;
			1407: d = 0;
			1408: d = 0;
			1409: d = 0;
			1410: d = 0;
			1411: d = 0;
			1412: d = 1;
			1413: d = 1;
			1414: d = 0;
			1415: d = 1;
			1416: d = 1;
			1417: d = 0;
			1418: d = 0;
			1419: d = 1;
			1420: d = 1;
			1421: d = 1;
			1422: d = 0;
			1423: d = 0;
			1424: d = 0;
			1425: d = 0;
			1426: d = 0;
			1427: d = 0;
			1428: d = 0;
			1429: d = 1;
			1430: d = 0;
			1431: d = 0;
			1432: d = 0;
			1433: d = 0;
			1434: d = 0;
			1435: d = 0;
			1436: d = 0;
			1437: d = 0;
			1438: d = 0;
			1439: d = 0;
			1440: d = 0;
			1441: d = 0;
			1442: d = 0;
			1443: d = 0;
			1444: d = 0;
			1445: d = 0;
			1446: d = 0;
			1447: d = 0;
			1448: d = 1;
			1449: d = 1;
			1450: d = 1;
			1451: d = 0;
			1452: d = 0;
			1453: d = 1;
			1454: d = 0;
			1455: d = 0;
			1456: d = 0;
			1457: d = 0;
			1458: d = 0;
			1459: d = 0;
			1460: d = 0;
			1461: d = 0;
			1462: d = 1;
			1463: d = 1;
			1464: d = 0;
			1465: d = 0;
			1466: d = 0;
			1467: d = 0;
			1468: d = 0;
			1469: d = 0;
			1470: d = 0;
			1471: d = 0;
			1472: d = 0;
			1473: d = 0;
			1474: d = 0;
			1475: d = 0;
			1476: d = 0;
			1477: d = 0;
			1478: d = 0;
			1479: d = 0;
			1480: d = 1;
			1481: d = 0;
			1482: d = 0;
			1483: d = 1;
			1484: d = 1;
			1485: d = 1;
			1486: d = 0;
			1487: d = 1;
			1488: d = 0;
			1489: d = 0;
			1490: d = 0;
			1491: d = 0;
			1492: d = 0;
			1493: d = 0;
			1494: d = 1;
			1495: d = 1;
			1496: d = 0;
			1497: d = 0;
			1498: d = 0;
			1499: d = 0;
			1500: d = 0;
			1501: d = 0;
			1502: d = 0;
			1503: d = 0;
			1504: d = 0;
			1505: d = 0;
			1506: d = 0;
			1507: d = 0;
			1508: d = 0;
			1509: d = 0;
			1510: d = 0;
			1511: d = 0;
			1512: d = 0;
			1513: d = 0;
			1514: d = 1;
			1515: d = 0;
			1516: d = 0;
			1517: d = 1;
			1518: d = 1;
			1519: d = 0;
			1520: d = 0;
			1521: d = 0;
			1522: d = 0;
			1523: d = 0;
			1524: d = 0;
			1525: d = 0;
			1526: d = 1;
			1527: d = 1;
			1528: d = 0;
			1529: d = 0;
			1530: d = 0;
			1531: d = 0;
			1532: d = 0;
			1533: d = 0;
			1534: d = 0;
			1535: d = 0;
			1536: d = 0;
			1537: d = 0;
			1538: d = 0;
			1539: d = 0;
			1540: d = 0;
			1541: d = 0;
			1542: d = 1;
			1543: d = 0;
			1544: d = 0;
			1545: d = 1;
			1546: d = 1;
			1547: d = 0;
			1548: d = 0;
			1549: d = 1;
			1550: d = 0;
			1551: d = 0;
			1552: d = 0;
			1553: d = 0;
			1554: d = 0;
			1555: d = 0;
			1556: d = 1;
			1557: d = 0;
			1558: d = 1;
			1559: d = 1;
			1560: d = 1;
			1561: d = 1;
			1562: d = 1;
			1563: d = 1;
			1564: d = 0;
			1565: d = 1;
			1566: d = 0;
			1567: d = 0;
			1568: d = 0;
			1569: d = 0;
			1570: d = 0;
			1571: d = 0;
			1572: d = 0;
			1573: d = 0;
			1574: d = 0;
			1575: d = 0;
			1576: d = 1;
			1577: d = 1;
			1578: d = 0;
			1579: d = 1;
			1580: d = 0;
			1581: d = 0;
			1582: d = 0;
			1583: d = 0;
			1584: d = 0;
			1585: d = 0;
			1586: d = 0;
			1587: d = 0;
			1588: d = 0;
			1589: d = 0;
			1590: d = 0;
			1591: d = 1;
			1592: d = 1;
			1593: d = 0;
			1594: d = 1;
			1595: d = 1;
			1596: d = 0;
			1597: d = 0;
			1598: d = 0;
			1599: d = 0;
			1600: d = 0;
			1601: d = 0;
			1602: d = 0;
			1603: d = 0;
			1604: d = 0;
			1605: d = 0;
			1606: d = 0;
			1607: d = 0;
			1608: d = 1;
			1609: d = 1;
			1610: d = 1;
			1611: d = 0;
			1612: d = 0;
			1613: d = 1;
			1614: d = 0;
			1615: d = 0;
			1616: d = 0;
			1617: d = 0;
			1618: d = 0;
			1619: d = 0;
			1620: d = 0;
			1621: d = 0;
			1622: d = 0;
			1623: d = 1;
			1624: d = 1;
			1625: d = 0;
			1626: d = 1;
			1627: d = 1;
			1628: d = 0;
			1629: d = 0;
			1630: d = 0;
			1631: d = 0;
			1632: d = 0;
			1633: d = 0;
			1634: d = 0;
			1635: d = 0;
			1636: d = 0;
			1637: d = 0;
			1638: d = 0;
			1639: d = 0;
			1640: d = 0;
			1641: d = 0;
			1642: d = 0;
			1643: d = 1;
			1644: d = 0;
			1645: d = 0;
			1646: d = 1;
			1647: d = 1;
			1648: d = 0;
			1649: d = 0;
			1650: d = 0;
			1651: d = 0;
			1652: d = 0;
			1653: d = 0;
			1654: d = 0;
			1655: d = 1;
			1656: d = 1;
			1657: d = 0;
			1658: d = 1;
			1659: d = 1;
			1660: d = 0;
			1661: d = 0;
			1662: d = 0;
			1663: d = 0;
			1664: d = 0;
			1665: d = 0;
			1666: d = 0;
			1667: d = 0;
			1668: d = 1;
			1669: d = 0;
			1670: d = 0;
			1671: d = 1;
			1672: d = 1;
			1673: d = 0;
			1674: d = 0;
			1675: d = 1;
			1676: d = 1;
			1677: d = 0;
			1678: d = 0;
			1679: d = 0;
			1680: d = 0;
			1681: d = 0;
			1682: d = 0;
			1683: d = 0;
			1684: d = 1;
			1685: d = 1;
			1686: d = 0;
			1687: d = 0;
			1688: d = 1;
			1689: d = 0;
			1690: d = 0;
			1691: d = 1;
			1692: d = 0;
			1693: d = 0;
			1694: d = 0;
			1695: d = 0;
			1696: d = 0;
			1697: d = 0;
			1698: d = 0;
			1699: d = 0;
			1700: d = 0;
			1701: d = 0;
			1702: d = 0;
			1703: d = 0;
			1704: d = 0;
			1705: d = 0;
			1706: d = 1;
			1707: d = 0;
			1708: d = 1;
			1709: d = 1;
			1710: d = 0;
			1711: d = 0;
			1712: d = 0;
			1713: d = 0;
			1714: d = 0;
			1715: d = 0;
			1716: d = 0;
			1717: d = 0;
			1718: d = 1;
			1719: d = 0;
			1720: d = 0;
			1721: d = 1;
			1722: d = 1;
			1723: d = 1;
			1724: d = 0;
			1725: d = 0;
			1726: d = 0;
			1727: d = 0;
			1728: d = 0;
			1729: d = 0;
			1730: d = 0;
			1731: d = 0;
			1732: d = 0;
			1733: d = 0;
			1734: d = 0;
			1735: d = 0;
			1736: d = 1;
			1737: d = 1;
			1738: d = 0;
			1739: d = 1;
			1740: d = 1;
			1741: d = 0;
			1742: d = 0;
			1743: d = 0;
			1744: d = 0;
			1745: d = 0;
			1746: d = 0;
			1747: d = 0;
			1748: d = 0;
			1749: d = 0;
			1750: d = 1;
			1751: d = 0;
			1752: d = 0;
			1753: d = 1;
			1754: d = 1;
			1755: d = 1;
			1756: d = 0;
			1757: d = 0;
			1758: d = 0;
			1759: d = 0;
			1760: d = 0;
			1761: d = 0;
			1762: d = 0;
			1763: d = 0;
			1764: d = 0;
			1765: d = 0;
			1766: d = 0;
			1767: d = 0;
			1768: d = 0;
			1769: d = 0;
			1770: d = 1;
			1771: d = 0;
			1772: d = 1;
			1773: d = 1;
			1774: d = 0;
			1775: d = 1;
			1776: d = 0;
			1777: d = 0;
			1778: d = 0;
			1779: d = 0;
			1780: d = 0;
			1781: d = 0;
			1782: d = 1;
			1783: d = 0;
			1784: d = 0;
			1785: d = 1;
			1786: d = 1;
			1787: d = 1;
			1788: d = 0;
			1789: d = 0;
			1790: d = 0;
			1791: d = 0;
			1792: d = 0;
			1793: d = 0;
			1794: d = 0;
			1795: d = 0;
			1796: d = 0;
			1797: d = 1;
			1798: d = 1;
			1799: d = 0;
			1800: d = 0;
			1801: d = 1;
			1802: d = 1;
			1803: d = 0;
			1804: d = 1;
			1805: d = 1;
			1806: d = 0;
			1807: d = 0;
			1808: d = 0;
			1809: d = 0;
			1810: d = 0;
			1811: d = 0;
			1812: d = 1;
			1813: d = 1;
			1814: d = 1;
			1815: d = 1;
			1816: d = 0;
			1817: d = 1;
			1818: d = 1;
			1819: d = 0;
			1820: d = 1;
			1821: d = 1;
			1822: d = 0;
			1823: d = 0;
			1824: d = 0;
			1825: d = 0;
			1826: d = 0;
			1827: d = 0;
			1828: d = 0;
			1829: d = 0;
			1830: d = 0;
			1831: d = 0;
			1832: d = 1;
			1833: d = 0;
			1834: d = 0;
			1835: d = 1;
			1836: d = 1;
			1837: d = 1;
			1838: d = 0;
			1839: d = 0;
			1840: d = 0;
			1841: d = 0;
			1842: d = 0;
			1843: d = 0;
			1844: d = 0;
			1845: d = 0;
			1846: d = 0;
			1847: d = 1;
			1848: d = 1;
			1849: d = 0;
			1850: d = 0;
			1851: d = 1;
			1852: d = 0;
			1853: d = 0;
			1854: d = 0;
			1855: d = 0;
			1856: d = 0;
			1857: d = 0;
			1858: d = 0;
			1859: d = 0;
			1860: d = 0;
			1861: d = 0;
			1862: d = 0;
			1863: d = 0;
			1864: d = 0;
			1865: d = 0;
			1866: d = 1;
			1867: d = 0;
			1868: d = 0;
			1869: d = 1;
			1870: d = 0;
			1871: d = 0;
			1872: d = 0;
			1873: d = 0;
			1874: d = 0;
			1875: d = 0;
			1876: d = 0;
			1877: d = 0;
			1878: d = 0;
			1879: d = 1;
			1880: d = 1;
			1881: d = 0;
			1882: d = 0;
			1883: d = 1;
			1884: d = 0;
			1885: d = 0;
			1886: d = 0;
			1887: d = 0;
			1888: d = 0;
			1889: d = 0;
			1890: d = 0;
			1891: d = 0;
			1892: d = 0;
			1893: d = 0;
			1894: d = 0;
			1895: d = 0;
			1896: d = 0;
			1897: d = 0;
			1898: d = 1;
			1899: d = 1;
			1900: d = 0;
			1901: d = 0;
			1902: d = 1;
			1903: d = 0;
			1904: d = 0;
			1905: d = 0;
			1906: d = 0;
			1907: d = 0;
			1908: d = 0;
			1909: d = 0;
			1910: d = 0;
			1911: d = 1;
			1912: d = 1;
			1913: d = 0;
			1914: d = 0;
			1915: d = 1;
			1916: d = 0;
			1917: d = 0;
			1918: d = 0;
			1919: d = 0;
			1920: d = 0;
			1921: d = 0;
			1922: d = 0;
			1923: d = 0;
			1924: d = 1;
			1925: d = 0;
			1926: d = 0;
			1927: d = 1;
			1928: d = 1;
			1929: d = 0;
			1930: d = 0;
			1931: d = 1;
			1932: d = 0;
			1933: d = 1;
			1934: d = 0;
			1935: d = 0;
			1936: d = 0;
			1937: d = 0;
			1938: d = 0;
			1939: d = 0;
			1940: d = 1;
			1941: d = 1;
			1942: d = 0;
			1943: d = 1;
			1944: d = 1;
			1945: d = 0;
			1946: d = 0;
			1947: d = 1;
			1948: d = 1;
			1949: d = 1;
			1950: d = 0;
			1951: d = 0;
			1952: d = 0;
			1953: d = 0;
			1954: d = 0;
			1955: d = 0;
			1956: d = 0;
			1957: d = 0;
			1958: d = 0;
			1959: d = 0;
			1960: d = 1;
			1961: d = 1;
			1962: d = 1;
			1963: d = 0;
			1964: d = 0;
			1965: d = 1;
			1966: d = 0;
			1967: d = 0;
			1968: d = 0;
			1969: d = 0;
			1970: d = 0;
			1971: d = 0;
			1972: d = 0;
			1973: d = 0;
			1974: d = 1;
			1975: d = 0;
			1976: d = 0;
			1977: d = 1;
			1978: d = 0;
			1979: d = 0;
			1980: d = 0;
			1981: d = 0;
			1982: d = 0;
			1983: d = 0;
			1984: d = 0;
			1985: d = 0;
			1986: d = 0;
			1987: d = 0;
			1988: d = 0;
			1989: d = 0;
			1990: d = 0;
			1991: d = 0;
			1992: d = 1;
			1993: d = 1;
			1994: d = 0;
			1995: d = 1;
			1996: d = 0;
			1997: d = 0;
			1998: d = 0;
			1999: d = 0;
			2000: d = 0;
			2001: d = 0;
			2002: d = 0;
			2003: d = 0;
			2004: d = 0;
			2005: d = 0;
			2006: d = 1;
			2007: d = 0;
			2008: d = 0;
			2009: d = 1;
			2010: d = 0;
			2011: d = 0;
			2012: d = 0;
			2013: d = 0;
			2014: d = 0;
			2015: d = 0;
			2016: d = 0;
			2017: d = 0;
			2018: d = 0;
			2019: d = 0;
			2020: d = 0;
			2021: d = 0;
			2022: d = 0;
			2023: d = 0;
			2024: d = 0;
			2025: d = 0;
			2026: d = 0;
			2027: d = 1;
			2028: d = 1;
			2029: d = 0;
			2030: d = 0;
			2031: d = 1;
			2032: d = 0;
			2033: d = 0;
			2034: d = 0;
			2035: d = 0;
			2036: d = 0;
			2037: d = 0;
			2038: d = 1;
			2039: d = 0;
			2040: d = 0;
			2041: d = 1;
			2042: d = 0;
			2043: d = 0;
			2044: d = 0;
			2045: d = 0;
			2046: d = 0;
			2047: d = 0;
			2048: d = 0;
			2049: d = 0;
			2050: d = 0;
			2051: d = 0;
			2052: d = 0;
			2053: d = 1;
			2054: d = 1;
			2055: d = 0;
			2056: d = 1;
			2057: d = 1;
			2058: d = 0;
			2059: d = 0;
			2060: d = 1;
			2061: d = 0;
			2062: d = 0;
			2063: d = 0;
			2064: d = 0;
			2065: d = 0;
			2066: d = 0;
			2067: d = 0;
			2068: d = 0;
			2069: d = 0;
			2070: d = 1;
			2071: d = 0;
			2072: d = 0;
			2073: d = 1;
			2074: d = 1;
			2075: d = 0;
			2076: d = 0;
			2077: d = 1;
			2078: d = 0;
			2079: d = 0;
			2080: d = 0;
			2081: d = 0;
			2082: d = 0;
			2083: d = 0;
			2084: d = 0;
			2085: d = 0;
			2086: d = 0;
			2087: d = 0;
			2088: d = 1;
			2089: d = 1;
			2090: d = 0;
			2091: d = 1;
			2092: d = 1;
			2093: d = 0;
			2094: d = 0;
			2095: d = 0;
			2096: d = 0;
			2097: d = 0;
			2098: d = 0;
			2099: d = 0;
			2100: d = 0;
			2101: d = 0;
			2102: d = 0;
			2103: d = 1;
			2104: d = 1;
			2105: d = 0;
			2106: d = 0;
			2107: d = 1;
			2108: d = 0;
			2109: d = 0;
			2110: d = 0;
			2111: d = 0;
			2112: d = 0;
			2113: d = 0;
			2114: d = 0;
			2115: d = 0;
			2116: d = 0;
			2117: d = 0;
			2118: d = 1;
			2119: d = 0;
			2120: d = 1;
			2121: d = 1;
			2122: d = 0;
			2123: d = 0;
			2124: d = 1;
			2125: d = 0;
			2126: d = 0;
			2127: d = 0;
			2128: d = 0;
			2129: d = 0;
			2130: d = 0;
			2131: d = 0;
			2132: d = 0;
			2133: d = 0;
			2134: d = 0;
			2135: d = 1;
			2136: d = 1;
			2137: d = 0;
			2138: d = 0;
			2139: d = 1;
			2140: d = 0;
			2141: d = 0;
			2142: d = 0;
			2143: d = 0;
			2144: d = 0;
			2145: d = 0;
			2146: d = 0;
			2147: d = 0;
			2148: d = 0;
			2149: d = 0;
			2150: d = 0;
			2151: d = 0;
			2152: d = 0;
			2153: d = 0;
			2154: d = 0;
			2155: d = 0;
			2156: d = 0;
			2157: d = 1;
			2158: d = 0;
			2159: d = 0;
			2160: d = 0;
			2161: d = 0;
			2162: d = 0;
			2163: d = 0;
			2164: d = 0;
			2165: d = 0;
			2166: d = 0;
			2167: d = 1;
			2168: d = 1;
			2169: d = 0;
			2170: d = 0;
			2171: d = 1;
			2172: d = 0;
			2173: d = 0;
			2174: d = 0;
			2175: d = 0;
			2176: d = 0;
			2177: d = 0;
			2178: d = 0;
			2179: d = 0;
			2180: d = 1;
			2181: d = 0;
			2182: d = 0;
			2183: d = 1;
			2184: d = 0;
			2185: d = 1;
			2186: d = 1;
			2187: d = 0;
			2188: d = 0;
			2189: d = 1;
			2190: d = 0;
			2191: d = 0;
			2192: d = 0;
			2193: d = 0;
			2194: d = 0;
			2195: d = 0;
			2196: d = 1;
			2197: d = 0;
			2198: d = 0;
			2199: d = 1;
			2200: d = 1;
			2201: d = 0;
			2202: d = 0;
			2203: d = 1;
			2204: d = 0;
			2205: d = 0;
			2206: d = 0;
			2207: d = 0;
			2208: d = 0;
			2209: d = 0;
			2210: d = 0;
			2211: d = 0;
			2212: d = 0;
			2213: d = 0;
			2214: d = 1;
			2215: d = 0;
			2216: d = 0;
			2217: d = 1;
			2218: d = 1;
			2219: d = 0;
			2220: d = 1;
			2221: d = 1;
			2222: d = 0;
			2223: d = 0;
			2224: d = 0;
			2225: d = 0;
			2226: d = 0;
			2227: d = 0;
			2228: d = 0;
			2229: d = 0;
			2230: d = 1;
			2231: d = 0;
			2232: d = 0;
			2233: d = 1;
			2234: d = 0;
			2235: d = 0;
			2236: d = 0;
			2237: d = 0;
			2238: d = 0;
			2239: d = 0;
			2240: d = 0;
			2241: d = 0;
			2242: d = 0;
			2243: d = 0;
			2244: d = 1;
			2245: d = 0;
			2246: d = 0;
			2247: d = 1;
			2248: d = 0;
			2249: d = 1;
			2250: d = 1;
			2251: d = 0;
			2252: d = 0;
			2253: d = 1;
			2254: d = 0;
			2255: d = 0;
			2256: d = 0;
			2257: d = 0;
			2258: d = 0;
			2259: d = 0;
			2260: d = 0;
			2261: d = 0;
			2262: d = 1;
			2263: d = 0;
			2264: d = 0;
			2265: d = 1;
			2266: d = 0;
			2267: d = 0;
			2268: d = 0;
			2269: d = 0;
			2270: d = 0;
			2271: d = 0;
			2272: d = 0;
			2273: d = 0;
			2274: d = 0;
			2275: d = 0;
			2276: d = 0;
			2277: d = 0;
			2278: d = 0;
			2279: d = 0;
			2280: d = 1;
			2281: d = 0;
			2282: d = 0;
			2283: d = 0;
			2284: d = 1;
			2285: d = 0;
			2286: d = 1;
			2287: d = 1;
			2288: d = 0;
			2289: d = 0;
			2290: d = 0;
			2291: d = 0;
			2292: d = 0;
			2293: d = 0;
			2294: d = 1;
			2295: d = 0;
			2296: d = 0;
			2297: d = 1;
			2298: d = 0;
			2299: d = 0;
			2300: d = 0;
			2301: d = 0;
			2302: d = 0;
			2303: d = 0;
			2304: d = 0;
			2305: d = 0;
			2306: d = 0;
			2307: d = 0;
			2308: d = 1;
			2309: d = 1;
			2310: d = 0;
			2311: d = 0;
			2312: d = 1;
			2313: d = 0;
			2314: d = 0;
			2315: d = 1;
			2316: d = 0;
			2317: d = 0;
			2318: d = 0;
			2319: d = 0;
			2320: d = 0;
			2321: d = 0;
			2322: d = 0;
			2323: d = 0;
			2324: d = 1;
			2325: d = 1;
			2326: d = 1;
			2327: d = 1;
			2328: d = 0;
			2329: d = 1;
			2330: d = 1;
			2331: d = 0;
			2332: d = 1;
			2333: d = 1;
			2334: d = 0;
			2335: d = 0;
			2336: d = 0;
			2337: d = 0;
			2338: d = 0;
			2339: d = 0;
			2340: d = 0;
			2341: d = 0;
			2342: d = 0;
			2343: d = 1;
			2344: d = 1;
			2345: d = 0;
			2346: d = 1;
			2347: d = 1;
			2348: d = 0;
			2349: d = 0;
			2350: d = 0;
			2351: d = 0;
			2352: d = 0;
			2353: d = 0;
			2354: d = 0;
			2355: d = 0;
			2356: d = 0;
			2357: d = 0;
			2358: d = 1;
			2359: d = 1;
			2360: d = 0;
			2361: d = 0;
			2362: d = 0;
			2363: d = 0;
			2364: d = 0;
			2365: d = 0;
			2366: d = 0;
			2367: d = 0;
			2368: d = 0;
			2369: d = 0;
			2370: d = 0;
			2371: d = 0;
			2372: d = 1;
			2373: d = 1;
			2374: d = 0;
			2375: d = 0;
			2376: d = 1;
			2377: d = 1;
			2378: d = 1;
			2379: d = 1;
			2380: d = 1;
			2381: d = 1;
			2382: d = 0;
			2383: d = 0;
			2384: d = 0;
			2385: d = 0;
			2386: d = 0;
			2387: d = 0;
			2388: d = 0;
			2389: d = 0;
			2390: d = 1;
			2391: d = 1;
			2392: d = 0;
			2393: d = 0;
			2394: d = 0;
			2395: d = 0;
			2396: d = 0;
			2397: d = 0;
			2398: d = 0;
			2399: d = 0;
			2400: d = 0;
			2401: d = 0;
			2402: d = 0;
			2403: d = 0;
			2404: d = 0;
			2405: d = 0;
			2406: d = 0;
			2407: d = 0;
			2408: d = 0;
			2409: d = 1;
			2410: d = 1;
			2411: d = 0;
			2412: d = 0;
			2413: d = 1;
			2414: d = 0;
			2415: d = 1;
			2416: d = 0;
			2417: d = 0;
			2418: d = 0;
			2419: d = 0;
			2420: d = 0;
			2421: d = 0;
			2422: d = 1;
			2423: d = 1;
			2424: d = 0;
			2425: d = 0;
			2426: d = 0;
			2427: d = 0;
			2428: d = 0;
			2429: d = 0;
			2430: d = 0;
			2431: d = 0;
			2432: d = 0;
			2433: d = 0;
			2434: d = 0;
			2435: d = 0;
			2436: d = 1;
			2437: d = 1;
			2438: d = 1;
			2439: d = 0;
			2440: d = 1;
			2441: d = 1;
			2442: d = 1;
			2443: d = 1;
			2444: d = 0;
			2445: d = 1;
			2446: d = 0;
			2447: d = 0;
			2448: d = 0;
			2449: d = 0;
			2450: d = 0;
			2451: d = 0;
			2452: d = 1;
			2453: d = 1;
			2454: d = 0;
			2455: d = 1;
			2456: d = 1;
			2457: d = 0;
			2458: d = 0;
			2459: d = 1;
			2460: d = 1;
			2461: d = 1;
			2462: d = 0;
			2463: d = 0;
			2464: d = 0;
			2465: d = 0;
			2466: d = 0;
			2467: d = 0;
			2468: d = 0;
			2469: d = 0;
			2470: d = 0;
			2471: d = 0;
			2472: d = 1;
			2473: d = 1;
			2474: d = 0;
			2475: d = 0;
			2476: d = 0;
			2477: d = 0;
			2478: d = 0;
			2479: d = 0;
			2480: d = 0;
			2481: d = 0;
			2482: d = 0;
			2483: d = 0;
			2484: d = 0;
			2485: d = 0;
			2486: d = 0;
			2487: d = 1;
			2488: d = 1;
			2489: d = 0;
			2490: d = 1;
			2491: d = 1;
			2492: d = 0;
			2493: d = 0;
			2494: d = 1;
			2495: d = 0;
			2496: d = 0;
			2497: d = 0;
			2498: d = 0;
			2499: d = 0;
			2500: d = 0;
			2501: d = 1;
			2502: d = 0;
			2503: d = 0;
			2504: d = 0;
			2505: d = 1;
			2506: d = 0;
			2507: d = 0;
			2508: d = 0;
			2509: d = 0;
			2510: d = 0;
			2511: d = 0;
			2512: d = 0;
			2513: d = 0;
			2514: d = 0;
			2515: d = 0;
			2516: d = 0;
			2517: d = 0;
			2518: d = 0;
			2519: d = 1;
			2520: d = 1;
			2521: d = 0;
			2522: d = 1;
			2523: d = 1;
			2524: d = 0;
			2525: d = 0;
			2526: d = 1;
			2527: d = 0;
			2528: d = 0;
			2529: d = 0;
			2530: d = 0;
			2531: d = 0;
			2532: d = 0;
			2533: d = 0;
			2534: d = 0;
			2535: d = 0;
			2536: d = 0;
			2537: d = 0;
			2538: d = 1;
			2539: d = 1;
			2540: d = 0;
			2541: d = 0;
			2542: d = 0;
			2543: d = 0;
			2544: d = 0;
			2545: d = 0;
			2546: d = 0;
			2547: d = 0;
			2548: d = 0;
			2549: d = 0;
			2550: d = 0;
			2551: d = 1;
			2552: d = 1;
			2553: d = 0;
			2554: d = 1;
			2555: d = 1;
			2556: d = 0;
			2557: d = 0;
			2558: d = 1;
			2559: d = 0;
			2560: d = 0;
			2561: d = 0;
			2562: d = 0;
			2563: d = 0;
			2564: d = 0;
			2565: d = 1;
			2566: d = 0;
			2567: d = 0;
			2568: d = 1;
			2569: d = 0;
			2570: d = 0;
			2571: d = 1;
			2572: d = 1;
			2573: d = 0;
			2574: d = 0;
			2575: d = 0;
			2576: d = 0;
			2577: d = 0;
			2578: d = 0;
			2579: d = 0;
			2580: d = 0;
			2581: d = 0;
			2582: d = 1;
			2583: d = 0;
			2584: d = 0;
			2585: d = 1;
			2586: d = 1;
			2587: d = 0;
			2588: d = 1;
			2589: d = 1;
			2590: d = 0;
			2591: d = 0;
			2592: d = 0;
			2593: d = 0;
			2594: d = 0;
			2595: d = 0;
			2596: d = 0;
			2597: d = 0;
			2598: d = 0;
			2599: d = 0;
			2600: d = 0;
			2601: d = 1;
			2602: d = 0;
			2603: d = 0;
			2604: d = 1;
			2605: d = 0;
			2606: d = 0;
			2607: d = 0;
			2608: d = 0;
			2609: d = 0;
			2610: d = 0;
			2611: d = 0;
			2612: d = 0;
			2613: d = 0;
			2614: d = 1;
			2615: d = 0;
			2616: d = 0;
			2617: d = 1;
			2618: d = 0;
			2619: d = 1;
			2620: d = 0;
			2621: d = 0;
			2622: d = 1;
			2623: d = 1;
			2624: d = 0;
			2625: d = 0;
			2626: d = 0;
			2627: d = 0;
			2628: d = 0;
			2629: d = 0;
			2630: d = 0;
			2631: d = 0;
			2632: d = 0;
			2633: d = 0;
			2634: d = 0;
			2635: d = 0;
			2636: d = 1;
			2637: d = 0;
			2638: d = 0;
			2639: d = 0;
			2640: d = 0;
			2641: d = 0;
			2642: d = 0;
			2643: d = 0;
			2644: d = 0;
			2645: d = 0;
			2646: d = 1;
			2647: d = 0;
			2648: d = 0;
			2649: d = 1;
			2650: d = 0;
			2651: d = 1;
			2652: d = 0;
			2653: d = 0;
			2654: d = 1;
			2655: d = 1;
			2656: d = 0;
			2657: d = 0;
			2658: d = 0;
			2659: d = 0;
			2660: d = 0;
			2661: d = 0;
			2662: d = 0;
			2663: d = 0;
			2664: d = 0;
			2665: d = 0;
			2666: d = 0;
			2667: d = 1;
			2668: d = 0;
			2669: d = 0;
			2670: d = 1;
			2671: d = 0;
			2672: d = 0;
			2673: d = 0;
			2674: d = 0;
			2675: d = 0;
			2676: d = 0;
			2677: d = 0;
			2678: d = 1;
			2679: d = 0;
			2680: d = 0;
			2681: d = 1;
			2682: d = 0;
			2683: d = 1;
			2684: d = 0;
			2685: d = 0;
			2686: d = 1;
			2687: d = 1;
			2688: d = 0;
			2689: d = 0;
			2690: d = 0;
			2691: d = 0;
			2692: d = 1;
			2693: d = 0;
			2694: d = 1;
			2695: d = 0;
			2696: d = 0;
			2697: d = 1;
			2698: d = 1;
			2699: d = 0;
			2700: d = 0;
			2701: d = 1;
			2702: d = 0;
			2703: d = 0;
			2704: d = 0;
			2705: d = 0;
			2706: d = 0;
			2707: d = 0;
			2708: d = 1;
			2709: d = 0;
			2710: d = 0;
			2711: d = 1;
			2712: d = 1;
			2713: d = 0;
			2714: d = 0;
			2715: d = 1;
			2716: d = 1;
			2717: d = 1;
			2718: d = 0;
			2719: d = 0;
			2720: d = 0;
			2721: d = 0;
			2722: d = 0;
			2723: d = 0;
			2724: d = 0;
			2725: d = 0;
			2726: d = 0;
			2727: d = 0;
			2728: d = 0;
			2729: d = 0;
			2730: d = 0;
			2731: d = 0;
			2732: d = 0;
			2733: d = 1;
			2734: d = 0;
			2735: d = 0;
			2736: d = 0;
			2737: d = 0;
			2738: d = 0;
			2739: d = 0;
			2740: d = 1;
			2741: d = 0;
			2742: d = 0;
			2743: d = 1;
			2744: d = 0;
			2745: d = 0;
			2746: d = 0;
			2747: d = 0;
			2748: d = 0;
			2749: d = 0;
			2750: d = 1;
			2751: d = 1;
			2752: d = 0;
			2753: d = 0;
			2754: d = 0;
			2755: d = 0;
			2756: d = 0;
			2757: d = 0;
			2758: d = 0;
			2759: d = 0;
			2760: d = 0;
			2761: d = 0;
			2762: d = 0;
			2763: d = 0;
			2764: d = 0;
			2765: d = 1;
			2766: d = 0;
			2767: d = 0;
			2768: d = 0;
			2769: d = 0;
			2770: d = 0;
			2771: d = 0;
			2772: d = 1;
			2773: d = 0;
			2774: d = 0;
			2775: d = 1;
			2776: d = 0;
			2777: d = 0;
			2778: d = 0;
			2779: d = 0;
			2780: d = 0;
			2781: d = 0;
			2782: d = 1;
			2783: d = 1;
			2784: d = 0;
			2785: d = 0;
			2786: d = 0;
			2787: d = 0;
			2788: d = 0;
			2789: d = 0;
			2790: d = 0;
			2791: d = 0;
			2792: d = 0;
			2793: d = 0;
			2794: d = 0;
			2795: d = 0;
			2796: d = 0;
			2797: d = 0;
			2798: d = 0;
			2799: d = 1;
			2800: d = 0;
			2801: d = 0;
			2802: d = 0;
			2803: d = 0;
			2804: d = 1;
			2805: d = 0;
			2806: d = 0;
			2807: d = 1;
			2808: d = 0;
			2809: d = 0;
			2810: d = 0;
			2811: d = 0;
			2812: d = 0;
			2813: d = 0;
			2814: d = 1;
			2815: d = 1;
			2816: d = 0;
			2817: d = 0;
			2818: d = 0;
			2819: d = 0;
			2820: d = 1;
			2821: d = 1;
			2822: d = 0;
			2823: d = 0;
			2824: d = 1;
			2825: d = 0;
			2826: d = 0;
			2827: d = 1;
			2828: d = 1;
			2829: d = 0;
			2830: d = 0;
			2831: d = 0;
			2832: d = 0;
			2833: d = 0;
			2834: d = 0;
			2835: d = 0;
			2836: d = 0;
			2837: d = 1;
			2838: d = 1;
			2839: d = 0;
			2840: d = 0;
			2841: d = 1;
			2842: d = 1;
			2843: d = 0;
			2844: d = 0;
			2845: d = 1;
			2846: d = 1;
			2847: d = 0;
			2848: d = 0;
			2849: d = 0;
			2850: d = 0;
			2851: d = 0;
			2852: d = 0;
			2853: d = 0;
			2854: d = 0;
			2855: d = 0;
			2856: d = 1;
			2857: d = 0;
			2858: d = 0;
			2859: d = 0;
			2860: d = 0;
			2861: d = 0;
			2862: d = 0;
			2863: d = 0;
			2864: d = 0;
			2865: d = 0;
			2866: d = 0;
			2867: d = 0;
			2868: d = 0;
			2869: d = 1;
			2870: d = 0;
			2871: d = 0;
			2872: d = 1;
			2873: d = 0;
			2874: d = 1;
			2875: d = 1;
			2876: d = 1;
			2877: d = 0;
			2878: d = 0;
			2879: d = 1;
			2880: d = 0;
			2881: d = 0;
			2882: d = 0;
			2883: d = 0;
			2884: d = 0;
			2885: d = 0;
			2886: d = 0;
			2887: d = 0;
			2888: d = 1;
			2889: d = 0;
			2890: d = 0;
			2891: d = 0;
			2892: d = 0;
			2893: d = 0;
			2894: d = 0;
			2895: d = 0;
			2896: d = 0;
			2897: d = 0;
			2898: d = 0;
			2899: d = 0;
			2900: d = 0;
			2901: d = 1;
			2902: d = 0;
			2903: d = 0;
			2904: d = 1;
			2905: d = 0;
			2906: d = 1;
			2907: d = 1;
			2908: d = 1;
			2909: d = 0;
			2910: d = 0;
			2911: d = 1;
			2912: d = 0;
			2913: d = 0;
			2914: d = 0;
			2915: d = 0;
			2916: d = 0;
			2917: d = 0;
			2918: d = 0;
			2919: d = 0;
			2920: d = 0;
			2921: d = 0;
			2922: d = 1;
			2923: d = 0;
			2924: d = 0;
			2925: d = 0;
			2926: d = 0;
			2927: d = 0;
			2928: d = 0;
			2929: d = 0;
			2930: d = 0;
			2931: d = 0;
			2932: d = 0;
			2933: d = 1;
			2934: d = 0;
			2935: d = 0;
			2936: d = 1;
			2937: d = 0;
			2938: d = 1;
			2939: d = 1;
			2940: d = 1;
			2941: d = 0;
			2942: d = 0;
			2943: d = 1;
			2944: d = 0;
			2945: d = 0;
			2946: d = 0;
			2947: d = 0;
			2948: d = 1;
			2949: d = 1;
			2950: d = 1;
			2951: d = 0;
			2952: d = 0;
			2953: d = 1;
			2954: d = 1;
			2955: d = 0;
			2956: d = 0;
			2957: d = 1;
			2958: d = 0;
			2959: d = 0;
			2960: d = 0;
			2961: d = 0;
			2962: d = 0;
			2963: d = 0;
			2964: d = 1;
			2965: d = 0;
			2966: d = 0;
			2967: d = 1;
			2968: d = 1;
			2969: d = 0;
			2970: d = 0;
			2971: d = 1;
			2972: d = 1;
			2973: d = 0;
			2974: d = 1;
			2975: d = 1;
			2976: d = 0;
			2977: d = 0;
			2978: d = 0;
			2979: d = 0;
			2980: d = 0;
			2981: d = 0;
			2982: d = 0;
			2983: d = 0;
			2984: d = 0;
			2985: d = 1;
			2986: d = 0;
			2987: d = 0;
			2988: d = 0;
			2989: d = 0;
			2990: d = 0;
			2991: d = 0;
			2992: d = 0;
			2993: d = 0;
			2994: d = 0;
			2995: d = 0;
			2996: d = 0;
			2997: d = 0;
			2998: d = 1;
			2999: d = 0;
			3000: d = 0;
			3001: d = 1;
			3002: d = 1;
			3003: d = 1;
			3004: d = 0;
			3005: d = 1;
			3006: d = 0;
			3007: d = 0;
			3008: d = 0;
			3009: d = 0;
			3010: d = 0;
			3011: d = 0;
			3012: d = 0;
			3013: d = 0;
			3014: d = 0;
			3015: d = 0;
			3016: d = 0;
			3017: d = 1;
			3018: d = 0;
			3019: d = 0;
			3020: d = 0;
			3021: d = 0;
			3022: d = 0;
			3023: d = 0;
			3024: d = 0;
			3025: d = 0;
			3026: d = 0;
			3027: d = 0;
			3028: d = 0;
			3029: d = 0;
			3030: d = 1;
			3031: d = 0;
			3032: d = 0;
			3033: d = 1;
			3034: d = 1;
			3035: d = 1;
			3036: d = 0;
			3037: d = 1;
			3038: d = 0;
			3039: d = 0;
			3040: d = 0;
			3041: d = 0;
			3042: d = 0;
			3043: d = 0;
			3044: d = 0;
			3045: d = 0;
			3046: d = 0;
			3047: d = 0;
			3048: d = 0;
			3049: d = 0;
			3050: d = 0;
			3051: d = 1;
			3052: d = 0;
			3053: d = 0;
			3054: d = 0;
			3055: d = 0;
			3056: d = 0;
			3057: d = 0;
			3058: d = 0;
			3059: d = 0;
			3060: d = 0;
			3061: d = 0;
			3062: d = 1;
			3063: d = 0;
			3064: d = 0;
			3065: d = 1;
			3066: d = 1;
			3067: d = 1;
			3068: d = 0;
			3069: d = 1;
			3070: d = 0;
			3071: d = 0;
			3072: d = 0;
			3073: d = 0;
			3074: d = 0;
			3075: d = 0;
			3076: d = 1;
			3077: d = 1;
			3078: d = 0;
			3079: d = 1;
			3080: d = 1;
			3081: d = 0;
			3082: d = 0;
			3083: d = 1;
			3084: d = 1;
			3085: d = 0;
			3086: d = 0;
			3087: d = 0;
			3088: d = 0;
			3089: d = 0;
			3090: d = 0;
			3091: d = 0;
			3092: d = 0;
			3093: d = 1;
			3094: d = 1;
			3095: d = 0;
			3096: d = 0;
			3097: d = 1;
			3098: d = 1;
			3099: d = 0;
			3100: d = 1;
			3101: d = 1;
			3102: d = 1;
			3103: d = 1;
			3104: d = 0;
			3105: d = 0;
			3106: d = 0;
			3107: d = 0;
			3108: d = 0;
			3109: d = 0;
			3110: d = 0;
			3111: d = 0;
			3112: d = 0;
			3113: d = 0;
			3114: d = 0;
			3115: d = 0;
			3116: d = 0;
			3117: d = 0;
			3118: d = 0;
			3119: d = 0;
			3120: d = 0;
			3121: d = 0;
			3122: d = 0;
			3123: d = 0;
			3124: d = 0;
			3125: d = 0;
			3126: d = 0;
			3127: d = 1;
			3128: d = 1;
			3129: d = 0;
			3130: d = 0;
			3131: d = 1;
			3132: d = 0;
			3133: d = 0;
			3134: d = 0;
			3135: d = 0;
			3136: d = 0;
			3137: d = 0;
			3138: d = 0;
			3139: d = 0;
			3140: d = 0;
			3141: d = 0;
			3142: d = 0;
			3143: d = 0;
			3144: d = 0;
			3145: d = 0;
			3146: d = 0;
			3147: d = 0;
			3148: d = 0;
			3149: d = 0;
			3150: d = 0;
			3151: d = 0;
			3152: d = 0;
			3153: d = 0;
			3154: d = 0;
			3155: d = 0;
			3156: d = 0;
			3157: d = 0;
			3158: d = 0;
			3159: d = 1;
			3160: d = 1;
			3161: d = 0;
			3162: d = 0;
			3163: d = 1;
			3164: d = 0;
			3165: d = 0;
			3166: d = 0;
			3167: d = 0;
			3168: d = 0;
			3169: d = 0;
			3170: d = 0;
			3171: d = 0;
			3172: d = 0;
			3173: d = 0;
			3174: d = 0;
			3175: d = 0;
			3176: d = 0;
			3177: d = 0;
			3178: d = 0;
			3179: d = 0;
			3180: d = 0;
			3181: d = 0;
			3182: d = 0;
			3183: d = 0;
			3184: d = 0;
			3185: d = 0;
			3186: d = 0;
			3187: d = 0;
			3188: d = 0;
			3189: d = 0;
			3190: d = 0;
			3191: d = 1;
			3192: d = 1;
			3193: d = 0;
			3194: d = 0;
			3195: d = 1;
			3196: d = 0;
			3197: d = 0;
			3198: d = 0;
			3199: d = 0;
			3200: d = 0;
			3201: d = 0;
			3202: d = 0;
			3203: d = 0;
			3204: d = 1;
			3205: d = 1;
			3206: d = 1;
			3207: d = 0;
			3208: d = 0;
			3209: d = 1;
			3210: d = 1;
			3211: d = 0;
			3212: d = 0;
			3213: d = 1;
			3214: d = 0;
			3215: d = 0;
			3216: d = 0;
			3217: d = 0;
			3218: d = 0;
			3219: d = 0;
			3220: d = 1;
			3221: d = 0;
			3222: d = 0;
			3223: d = 1;
			3224: d = 1;
			3225: d = 0;
			3226: d = 0;
			3227: d = 0;
			3228: d = 1;
			3229: d = 0;
			3230: d = 0;
			3231: d = 1;
			3232: d = 0;
			3233: d = 0;
			3234: d = 0;
			3235: d = 0;
			3236: d = 0;
			3237: d = 0;
			3238: d = 0;
			3239: d = 0;
			3240: d = 0;
			3241: d = 0;
			3242: d = 0;
			3243: d = 0;
			3244: d = 0;
			3245: d = 0;
			3246: d = 0;
			3247: d = 0;
			3248: d = 0;
			3249: d = 0;
			3250: d = 0;
			3251: d = 0;
			3252: d = 0;
			3253: d = 0;
			3254: d = 1;
			3255: d = 0;
			3256: d = 0;
			3257: d = 1;
			3258: d = 0;
			3259: d = 0;
			3260: d = 0;
			3261: d = 0;
			3262: d = 0;
			3263: d = 0;
			3264: d = 0;
			3265: d = 0;
			3266: d = 0;
			3267: d = 0;
			3268: d = 0;
			3269: d = 0;
			3270: d = 0;
			3271: d = 0;
			3272: d = 0;
			3273: d = 0;
			3274: d = 0;
			3275: d = 0;
			3276: d = 0;
			3277: d = 0;
			3278: d = 0;
			3279: d = 0;
			3280: d = 0;
			3281: d = 0;
			3282: d = 0;
			3283: d = 0;
			3284: d = 0;
			3285: d = 0;
			3286: d = 1;
			3287: d = 0;
			3288: d = 0;
			3289: d = 1;
			3290: d = 0;
			3291: d = 0;
			3292: d = 0;
			3293: d = 0;
			3294: d = 0;
			3295: d = 0;
			3296: d = 0;
			3297: d = 0;
			3298: d = 0;
			3299: d = 0;
			3300: d = 0;
			3301: d = 0;
			3302: d = 0;
			3303: d = 0;
			3304: d = 0;
			3305: d = 0;
			3306: d = 0;
			3307: d = 0;
			3308: d = 0;
			3309: d = 0;
			3310: d = 0;
			3311: d = 0;
			3312: d = 0;
			3313: d = 0;
			3314: d = 0;
			3315: d = 0;
			3316: d = 0;
			3317: d = 0;
			3318: d = 1;
			3319: d = 0;
			3320: d = 0;
			3321: d = 1;
			3322: d = 0;
			3323: d = 0;
			3324: d = 0;
			3325: d = 0;
			3326: d = 0;
			3327: d = 0;
			3328: d = 0;
			3329: d = 0;
			3330: d = 0;
			3331: d = 0;
			3332: d = 1;
			3333: d = 1;
			3334: d = 0;
			3335: d = 0;
			3336: d = 1;
			3337: d = 0;
			3338: d = 1;
			3339: d = 1;
			3340: d = 1;
			3341: d = 1;
			3342: d = 0;
			3343: d = 0;
			3344: d = 0;
			3345: d = 0;
			3346: d = 0;
			3347: d = 0;
			3348: d = 0;
			3349: d = 1;
			3350: d = 1;
			3351: d = 0;
			3352: d = 1;
			3353: d = 1;
			3354: d = 1;
			3355: d = 0;
			3356: d = 0;
			3357: d = 1;
			3358: d = 0;
			3359: d = 0;
			3360: d = 0;
			3361: d = 0;
			3362: d = 0;
			3363: d = 0;
			3364: d = 0;
			3365: d = 0;
			3366: d = 0;
			3367: d = 0;
			3368: d = 0;
			3369: d = 0;
			3370: d = 0;
			3371: d = 0;
			3372: d = 0;
			3373: d = 0;
			3374: d = 0;
			3375: d = 0;
			3376: d = 0;
			3377: d = 0;
			3378: d = 0;
			3379: d = 0;
			3380: d = 0;
			3381: d = 0;
			3382: d = 0;
			3383: d = 1;
			3384: d = 0;
			3385: d = 0;
			3386: d = 0;
			3387: d = 0;
			3388: d = 0;
			3389: d = 0;
			3390: d = 0;
			3391: d = 0;
			3392: d = 0;
			3393: d = 0;
			3394: d = 0;
			3395: d = 0;
			3396: d = 0;
			3397: d = 0;
			3398: d = 0;
			3399: d = 0;
			3400: d = 0;
			3401: d = 0;
			3402: d = 0;
			3403: d = 0;
			3404: d = 0;
			3405: d = 0;
			3406: d = 0;
			3407: d = 0;
			3408: d = 0;
			3409: d = 0;
			3410: d = 0;
			3411: d = 0;
			3412: d = 0;
			3413: d = 0;
			3414: d = 0;
			3415: d = 1;
			3416: d = 0;
			3417: d = 0;
			3418: d = 0;
			3419: d = 0;
			3420: d = 0;
			3421: d = 0;
			3422: d = 0;
			3423: d = 0;
			3424: d = 0;
			3425: d = 0;
			3426: d = 0;
			3427: d = 0;
			3428: d = 0;
			3429: d = 0;
			3430: d = 0;
			3431: d = 0;
			3432: d = 0;
			3433: d = 0;
			3434: d = 0;
			3435: d = 0;
			3436: d = 0;
			3437: d = 0;
			3438: d = 0;
			3439: d = 0;
			3440: d = 0;
			3441: d = 0;
			3442: d = 0;
			3443: d = 0;
			3444: d = 0;
			3445: d = 0;
			3446: d = 0;
			3447: d = 1;
			3448: d = 0;
			3449: d = 0;
			3450: d = 0;
			3451: d = 0;
			3452: d = 0;
			3453: d = 0;
			3454: d = 0;
			3455: d = 0;
			3456: d = 0;
			3457: d = 0;
			3458: d = 0;
			3459: d = 0;
			3460: d = 0;
			3461: d = 1;
			3462: d = 0;
			3463: d = 0;
			3464: d = 0;
			3465: d = 0;
			3466: d = 0;
			3467: d = 0;
			3468: d = 0;
			3469: d = 0;
			3470: d = 0;
			3471: d = 0;
			3472: d = 0;
			3473: d = 0;
			3474: d = 0;
			3475: d = 0;
			3476: d = 1;
			3477: d = 0;
			3478: d = 0;
			3479: d = 1;
			3480: d = 1;
			3481: d = 1;
			3482: d = 0;
			3483: d = 1;
			3484: d = 0;
			3485: d = 0;
			3486: d = 0;
			3487: d = 0;
			3488: d = 0;
			3489: d = 0;
			3490: d = 0;
			3491: d = 0;
			3492: d = 0;
			3493: d = 0;
			3494: d = 0;
			3495: d = 0;
			3496: d = 0;
			3497: d = 0;
			3498: d = 0;
			3499: d = 0;
			3500: d = 0;
			3501: d = 0;
			3502: d = 0;
			3503: d = 0;
			3504: d = 0;
			3505: d = 0;
			3506: d = 0;
			3507: d = 0;
			3508: d = 0;
			3509: d = 0;
			3510: d = 0;
			3511: d = 0;
			3512: d = 0;
			3513: d = 0;
			3514: d = 0;
			3515: d = 0;
			3516: d = 0;
			3517: d = 0;
			3518: d = 0;
			3519: d = 0;
			3520: d = 0;
			3521: d = 0;
			3522: d = 0;
			3523: d = 0;
			3524: d = 0;
			3525: d = 0;
			3526: d = 0;
			3527: d = 0;
			3528: d = 0;
			3529: d = 0;
			3530: d = 0;
			3531: d = 0;
			3532: d = 0;
			3533: d = 0;
			3534: d = 0;
			3535: d = 0;
			3536: d = 0;
			3537: d = 0;
			3538: d = 0;
			3539: d = 0;
			3540: d = 0;
			3541: d = 0;
			3542: d = 0;
			3543: d = 0;
			3544: d = 0;
			3545: d = 0;
			3546: d = 0;
			3547: d = 0;
			3548: d = 0;
			3549: d = 0;
			3550: d = 0;
			3551: d = 0;
			3552: d = 0;
			3553: d = 0;
			3554: d = 0;
			3555: d = 0;
			3556: d = 0;
			3557: d = 0;
			3558: d = 0;
			3559: d = 0;
			3560: d = 0;
			3561: d = 0;
			3562: d = 0;
			3563: d = 0;
			3564: d = 0;
			3565: d = 0;
			3566: d = 0;
			3567: d = 0;
			3568: d = 0;
			3569: d = 0;
			3570: d = 0;
			3571: d = 0;
			3572: d = 0;
			3573: d = 0;
			3574: d = 0;
			3575: d = 0;
			3576: d = 0;
			3577: d = 0;
			3578: d = 0;
			3579: d = 0;
			3580: d = 0;
			3581: d = 0;
			3582: d = 0;
			3583: d = 0;
			3584: d = 0;
			3585: d = 0;
			3586: d = 0;
			3587: d = 0;
			3588: d = 1;
			3589: d = 0;
			3590: d = 1;
			3591: d = 1;
			3592: d = 1;
			3593: d = 1;
			3594: d = 1;
			3595: d = 1;
			3596: d = 1;
			3597: d = 1;
			3598: d = 0;
			3599: d = 0;
			3600: d = 0;
			3601: d = 0;
			3602: d = 0;
			3603: d = 0;
			3604: d = 1;
			3605: d = 1;
			3606: d = 0;
			3607: d = 0;
			3608: d = 0;
			3609: d = 0;
			3610: d = 0;
			3611: d = 0;
			3612: d = 0;
			3613: d = 0;
			3614: d = 0;
			3615: d = 0;
			3616: d = 0;
			3617: d = 0;
			3618: d = 0;
			3619: d = 0;
			3620: d = 0;
			3621: d = 0;
			3622: d = 0;
			3623: d = 0;
			3624: d = 0;
			3625: d = 0;
			3626: d = 0;
			3627: d = 0;
			3628: d = 0;
			3629: d = 0;
			3630: d = 0;
			3631: d = 0;
			3632: d = 0;
			3633: d = 0;
			3634: d = 0;
			3635: d = 0;
			3636: d = 0;
			3637: d = 0;
			3638: d = 0;
			3639: d = 0;
			3640: d = 0;
			3641: d = 0;
			3642: d = 0;
			3643: d = 0;
			3644: d = 0;
			3645: d = 0;
			3646: d = 0;
			3647: d = 0;
			3648: d = 0;
			3649: d = 0;
			3650: d = 0;
			3651: d = 0;
			3652: d = 0;
			3653: d = 0;
			3654: d = 0;
			3655: d = 0;
			3656: d = 0;
			3657: d = 0;
			3658: d = 0;
			3659: d = 0;
			3660: d = 0;
			3661: d = 0;
			3662: d = 0;
			3663: d = 0;
			3664: d = 0;
			3665: d = 0;
			3666: d = 0;
			3667: d = 0;
			3668: d = 0;
			3669: d = 0;
			3670: d = 0;
			3671: d = 0;
			3672: d = 0;
			3673: d = 0;
			3674: d = 0;
			3675: d = 0;
			3676: d = 0;
			3677: d = 0;
			3678: d = 0;
			3679: d = 0;
			3680: d = 0;
			3681: d = 0;
			3682: d = 0;
			3683: d = 0;
			3684: d = 0;
			3685: d = 0;
			3686: d = 0;
			3687: d = 0;
			3688: d = 0;
			3689: d = 0;
			3690: d = 0;
			3691: d = 0;
			3692: d = 0;
			3693: d = 0;
			3694: d = 0;
			3695: d = 0;
			3696: d = 0;
			3697: d = 0;
			3698: d = 0;
			3699: d = 0;
			3700: d = 0;
			3701: d = 0;
			3702: d = 0;
			3703: d = 0;
			3704: d = 0;
			3705: d = 0;
			3706: d = 0;
			3707: d = 0;
			3708: d = 0;
			3709: d = 0;
			3710: d = 0;
			3711: d = 0;
			3712: d = 0;
			3713: d = 0;
			3714: d = 0;
			3715: d = 0;
			3716: d = 0;
			3717: d = 1;
			3718: d = 0;
			3719: d = 0;
			3720: d = 0;
			3721: d = 0;
			3722: d = 0;
			3723: d = 0;
			3724: d = 1;
			3725: d = 1;
			3726: d = 0;
			3727: d = 0;
			3728: d = 0;
			3729: d = 0;
			3730: d = 0;
			3731: d = 0;
			3732: d = 1;
			3733: d = 1;
			3734: d = 0;
			3735: d = 1;
			3736: d = 0;
			3737: d = 0;
			3738: d = 0;
			3739: d = 0;
			3740: d = 0;
			3741: d = 0;
			3742: d = 0;
			3743: d = 0;
			3744: d = 0;
			3745: d = 0;
			3746: d = 0;
			3747: d = 0;
			3748: d = 0;
			3749: d = 0;
			3750: d = 0;
			3751: d = 0;
			3752: d = 0;
			3753: d = 0;
			3754: d = 0;
			3755: d = 0;
			3756: d = 0;
			3757: d = 0;
			3758: d = 0;
			3759: d = 0;
			3760: d = 0;
			3761: d = 0;
			3762: d = 0;
			3763: d = 0;
			3764: d = 0;
			3765: d = 0;
			3766: d = 0;
			3767: d = 0;
			3768: d = 0;
			3769: d = 0;
			3770: d = 0;
			3771: d = 0;
			3772: d = 0;
			3773: d = 0;
			3774: d = 0;
			3775: d = 0;
			3776: d = 0;
			3777: d = 0;
			3778: d = 0;
			3779: d = 0;
			3780: d = 0;
			3781: d = 0;
			3782: d = 0;
			3783: d = 0;
			3784: d = 0;
			3785: d = 0;
			3786: d = 0;
			3787: d = 0;
			3788: d = 0;
			3789: d = 0;
			3790: d = 0;
			3791: d = 0;
			3792: d = 0;
			3793: d = 0;
			3794: d = 0;
			3795: d = 0;
			3796: d = 0;
			3797: d = 0;
			3798: d = 0;
			3799: d = 0;
			3800: d = 0;
			3801: d = 0;
			3802: d = 0;
			3803: d = 0;
			3804: d = 0;
			3805: d = 0;
			3806: d = 0;
			3807: d = 0;
			3808: d = 0;
			3809: d = 0;
			3810: d = 0;
			3811: d = 0;
			3812: d = 0;
			3813: d = 0;
			3814: d = 0;
			3815: d = 0;
			3816: d = 0;
			3817: d = 0;
			3818: d = 0;
			3819: d = 0;
			3820: d = 0;
			3821: d = 0;
			3822: d = 0;
			3823: d = 0;
			3824: d = 0;
			3825: d = 0;
			3826: d = 0;
			3827: d = 0;
			3828: d = 0;
			3829: d = 0;
			3830: d = 0;
			3831: d = 0;
			3832: d = 0;
			3833: d = 0;
			3834: d = 0;
			3835: d = 0;
			3836: d = 0;
			3837: d = 0;
			3838: d = 0;
			3839: d = 0;
			3840: d = 1'bX;
			3841: d = 1'bX;
			3842: d = 1'bX;
			3843: d = 1'bX;
			3844: d = 1'bX;
			3845: d = 1'bX;
			3846: d = 1'bX;
			3847: d = 1'bX;
			3848: d = 1'bX;
			3849: d = 1'bX;
			3850: d = 1'bX;
			3851: d = 1'bX;
			3852: d = 1'bX;
			3853: d = 1'bX;
			3854: d = 1'bX;
			3855: d = 1'bX;
			3856: d = 1'bX;
			3857: d = 1'bX;
			3858: d = 1'bX;
			3859: d = 1'bX;
			3860: d = 1'bX;
			3861: d = 1'bX;
			3862: d = 1'bX;
			3863: d = 1'bX;
			3864: d = 1'bX;
			3865: d = 1'bX;
			3866: d = 1'bX;
			3867: d = 1'bX;
			3868: d = 1'bX;
			3869: d = 1'bX;
			3870: d = 1'bX;
			3871: d = 1'bX;
			3872: d = 1'bX;
			3873: d = 1'bX;
			3874: d = 1'bX;
			3875: d = 1'bX;
			3876: d = 1'bX;
			3877: d = 1'bX;
			3878: d = 1'bX;
			3879: d = 1'bX;
			3880: d = 1'bX;
			3881: d = 1'bX;
			3882: d = 1'bX;
			3883: d = 1'bX;
			3884: d = 1'bX;
			3885: d = 1'bX;
			3886: d = 1'bX;
			3887: d = 1'bX;
			3888: d = 1'bX;
			3889: d = 1'bX;
			3890: d = 1'bX;
			3891: d = 1'bX;
			3892: d = 1'bX;
			3893: d = 1'bX;
			3894: d = 1'bX;
			3895: d = 1'bX;
			3896: d = 1'bX;
			3897: d = 1'bX;
			3898: d = 1'bX;
			3899: d = 1'bX;
			3900: d = 1'bX;
			3901: d = 1'bX;
			3902: d = 1'bX;
			3903: d = 1'bX;
			3904: d = 1'bX;
			3905: d = 1'bX;
			3906: d = 1'bX;
			3907: d = 1'bX;
			3908: d = 1'bX;
			3909: d = 1'bX;
			3910: d = 1'bX;
			3911: d = 1'bX;
			3912: d = 1'bX;
			3913: d = 1'bX;
			3914: d = 1'bX;
			3915: d = 1'bX;
			3916: d = 1'bX;
			3917: d = 1'bX;
			3918: d = 1'bX;
			3919: d = 1'bX;
			3920: d = 1'bX;
			3921: d = 1'bX;
			3922: d = 1'bX;
			3923: d = 1'bX;
			3924: d = 1'bX;
			3925: d = 1'bX;
			3926: d = 1'bX;
			3927: d = 1'bX;
			3928: d = 1'bX;
			3929: d = 1'bX;
			3930: d = 1'bX;
			3931: d = 1'bX;
			3932: d = 1'bX;
			3933: d = 1'bX;
			3934: d = 1'bX;
			3935: d = 1'bX;
			3936: d = 1'bX;
			3937: d = 1'bX;
			3938: d = 1'bX;
			3939: d = 1'bX;
			3940: d = 1'bX;
			3941: d = 1'bX;
			3942: d = 1'bX;
			3943: d = 1'bX;
			3944: d = 1'bX;
			3945: d = 1'bX;
			3946: d = 1'bX;
			3947: d = 1'bX;
			3948: d = 1'bX;
			3949: d = 1'bX;
			3950: d = 1'bX;
			3951: d = 1'bX;
			3952: d = 1'bX;
			3953: d = 1'bX;
			3954: d = 1'bX;
			3955: d = 1'bX;
			3956: d = 1'bX;
			3957: d = 1'bX;
			3958: d = 1'bX;
			3959: d = 1'bX;
			3960: d = 1'bX;
			3961: d = 1'bX;
			3962: d = 1'bX;
			3963: d = 1'bX;
			3964: d = 1'bX;
			3965: d = 1'bX;
			3966: d = 1'bX;
			3967: d = 1'bX;
			3968: d = 1'bX;
			3969: d = 1'bX;
			3970: d = 1'bX;
			3971: d = 1'bX;
			3972: d = 1'bX;
			3973: d = 1'bX;
			3974: d = 1'bX;
			3975: d = 1'bX;
			3976: d = 1'bX;
			3977: d = 1'bX;
			3978: d = 1'bX;
			3979: d = 1'bX;
			3980: d = 1'bX;
			3981: d = 1'bX;
			3982: d = 1'bX;
			3983: d = 1'bX;
			3984: d = 1'bX;
			3985: d = 1'bX;
			3986: d = 1'bX;
			3987: d = 1'bX;
			3988: d = 1'bX;
			3989: d = 1'bX;
			3990: d = 1'bX;
			3991: d = 1'bX;
			3992: d = 1'bX;
			3993: d = 1'bX;
			3994: d = 1'bX;
			3995: d = 1'bX;
			3996: d = 1'bX;
			3997: d = 1'bX;
			3998: d = 1'bX;
			3999: d = 1'bX;
			4000: d = 1'bX;
			4001: d = 1'bX;
			4002: d = 1'bX;
			4003: d = 1'bX;
			4004: d = 1'bX;
			4005: d = 1'bX;
			4006: d = 1'bX;
			4007: d = 1'bX;
			4008: d = 1'bX;
			4009: d = 1'bX;
			4010: d = 1'bX;
			4011: d = 1'bX;
			4012: d = 1'bX;
			4013: d = 1'bX;
			4014: d = 1'bX;
			4015: d = 1'bX;
			4016: d = 1'bX;
			4017: d = 1'bX;
			4018: d = 1'bX;
			4019: d = 1'bX;
			4020: d = 1'bX;
			4021: d = 1'bX;
			4022: d = 1'bX;
			4023: d = 1'bX;
			4024: d = 1'bX;
			4025: d = 1'bX;
			4026: d = 1'bX;
			4027: d = 1'bX;
			4028: d = 1'bX;
			4029: d = 1'bX;
			4030: d = 1'bX;
			4031: d = 1'bX;
			4032: d = 1'bX;
			4033: d = 1'bX;
			4034: d = 1'bX;
			4035: d = 1'bX;
			4036: d = 1'bX;
			4037: d = 1'bX;
			4038: d = 1'bX;
			4039: d = 1'bX;
			4040: d = 1'bX;
			4041: d = 1'bX;
			4042: d = 1'bX;
			4043: d = 1'bX;
			4044: d = 1'bX;
			4045: d = 1'bX;
			4046: d = 1'bX;
			4047: d = 1'bX;
			4048: d = 1'bX;
			4049: d = 1'bX;
			4050: d = 1'bX;
			4051: d = 1'bX;
			4052: d = 1'bX;
			4053: d = 1'bX;
			4054: d = 1'bX;
			4055: d = 1'bX;
			4056: d = 1'bX;
			4057: d = 1'bX;
			4058: d = 1'bX;
			4059: d = 1'bX;
			4060: d = 1'bX;
			4061: d = 1'bX;
			4062: d = 1'bX;
			4063: d = 1'bX;
			4064: d = 1'bX;
			4065: d = 1'bX;
			4066: d = 1'bX;
			4067: d = 1'bX;
			4068: d = 1'bX;
			4069: d = 1'bX;
			4070: d = 1'bX;
			4071: d = 1'bX;
			4072: d = 1'bX;
			4073: d = 1'bX;
			4074: d = 1'bX;
			4075: d = 1'bX;
			4076: d = 1'bX;
			4077: d = 1'bX;
			4078: d = 1'bX;
			4079: d = 1'bX;
			4080: d = 1'bX;
			4081: d = 1'bX;
			4082: d = 1'bX;
			4083: d = 1'bX;
			4084: d = 1'bX;
			4085: d = 1'bX;
			4086: d = 1'bX;
			4087: d = 1'bX;
			4088: d = 1'bX;
			4089: d = 1'bX;
			4090: d = 1'bX;
			4091: d = 1'bX;
			4092: d = 1'bX;
			4093: d = 1'bX;
			4094: d = 1'bX;
			4095: d = 1'bX;
			default: d = 'X;
		endcase
	end

	assign data = d;
endmodule : logo_table
